netcdf land_hgrid {
dimensions:
	stringlen = 255 ;
	nxp = 289 ;
	nyp = 181 ;
	nx = 288 ;
	ny = 180 ;
variables:
	char tile(stringlen) ;
		tile:standard_name = "grid_tile_spec" ;
		tile:tile_spec_version = "0.2" ;
		tile:geometry = "spherical" ;
		tile:discretization = "logically_rectangular" ;
		tile:conformal = "true" ;
	double x(nyp, nxp) ;
		x:standard_name = "geographic_longitude" ;
		x:units = "degree_east" ;
	double y(nyp, nxp) ;
		y:standard_name = "geographic_latitude" ;
		y:units = "degree_north" ;
	double dx(nyp, nx) ;
		dx:standard_name = "grid_edge_x_distance" ;
		dx:units = "meters" ;
	double dy(ny, nxp) ;
		dy:standard_name = "grid_edge_y_distance" ;
		dy:units = "meters" ;
	double angle_dx(nyp, nxp) ;
		angle_dx:standard_name = "grid_vertex_x_angle_WRT_geographic_east" ;
		angle_dx:units = "degrees_east" ;
	double area(ny, nx) ;
		area:standard_name = "grid_cell_area" ;
		area:units = "m2" ;
data:

 tile = "tile1" ;

 x =
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360,
  0, 1.25, 2.5, 3.75, 5, 6.25, 7.5, 8.75, 10, 11.25, 12.5, 13.75, 15, 16.25, 
    17.5, 18.75, 20, 21.25, 22.5, 23.75, 25, 26.25, 27.5, 28.75, 30, 31.25, 
    32.5, 33.75, 35, 36.25, 37.5, 38.75, 40, 41.25, 42.5, 43.75, 45, 46.25, 
    47.5, 48.75, 50, 51.25, 52.5, 53.75, 55, 56.25, 57.5, 58.75, 60, 61.25, 
    62.5, 63.75, 65, 66.25, 67.5, 68.75, 70, 71.25, 72.5, 73.75, 75, 76.25, 
    77.5, 78.75, 80, 81.25, 82.5, 83.75, 85, 86.25, 87.5, 88.75, 90, 91.25, 
    92.5, 93.75, 95, 96.25, 97.5, 98.75, 100, 101.25, 102.5, 103.75, 105, 
    106.25, 107.5, 108.75, 110, 111.25, 112.5, 113.75, 115, 116.25, 117.5, 
    118.75, 120, 121.25, 122.5, 123.75, 125, 126.25, 127.5, 128.75, 130, 
    131.25, 132.5, 133.75, 135, 136.25, 137.5, 138.75, 140, 141.25, 142.5, 
    143.75, 145, 146.25, 147.5, 148.75, 150, 151.25, 152.5, 153.75, 155, 
    156.25, 157.5, 158.75, 160, 161.25, 162.5, 163.75, 165, 166.25, 167.5, 
    168.75, 170, 171.25, 172.5, 173.75, 175, 176.25, 177.5, 178.75, 180, 
    181.25, 182.5, 183.75, 185, 186.25, 187.5, 188.75, 190, 191.25, 192.5, 
    193.75, 195, 196.25, 197.5, 198.75, 200, 201.25, 202.5, 203.75, 205, 
    206.25, 207.5, 208.75, 210, 211.25, 212.5, 213.75, 215, 216.25, 217.5, 
    218.75, 220, 221.25, 222.5, 223.75, 225, 226.25, 227.5, 228.75, 230, 
    231.25, 232.5, 233.75, 235, 236.25, 237.5, 238.75, 240, 241.25, 242.5, 
    243.75, 245, 246.25, 247.5, 248.75, 250, 251.25, 252.5, 253.75, 255, 
    256.25, 257.5, 258.75, 260, 261.25, 262.5, 263.75, 265, 266.25, 267.5, 
    268.75, 270, 271.25, 272.5, 273.75, 275, 276.25, 277.5, 278.75, 280, 
    281.25, 282.5, 283.75, 285, 286.25, 287.5, 288.75, 290, 291.25, 292.5, 
    293.75, 295, 296.25, 297.5, 298.75, 300, 301.25, 302.5, 303.75, 305, 
    306.25, 307.5, 308.75, 310, 311.25, 312.5, 313.75, 315, 316.25, 317.5, 
    318.75, 320, 321.25, 322.5, 323.75, 325, 326.25, 327.5, 328.75, 330, 
    331.25, 332.5, 333.75, 335, 336.25, 337.5, 338.75, 340, 341.25, 342.5, 
    343.75, 345, 346.25, 347.5, 348.75, 350, 351.25, 352.5, 353.75, 355, 
    356.25, 357.5, 358.75, 360 ;

 y =
  -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, -90, 
    -90, -90, -90, -90, -90, -90, -90, -90,
  -89.4943820224719, -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719, 
    -89.4943820224719, -89.4943820224719, -89.4943820224719,
  -88.9887640449438, -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438, 
    -88.9887640449438, -88.9887640449438, -88.9887640449438,
  -87.9775280898876, -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876, 
    -87.9775280898876, -87.9775280898876, -87.9775280898876,
  -86.9662921348315, -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315, 
    -86.9662921348315, -86.9662921348315, -86.9662921348315,
  -85.9550561797753, -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753, 
    -85.9550561797753, -85.9550561797753, -85.9550561797753,
  -84.9438202247191, -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191, 
    -84.9438202247191, -84.9438202247191, -84.9438202247191,
  -83.9325842696629, -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629, 
    -83.9325842696629, -83.9325842696629, -83.9325842696629,
  -82.9213483146067, -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067, 
    -82.9213483146067, -82.9213483146067, -82.9213483146067,
  -81.9101123595506, -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506, 
    -81.9101123595506, -81.9101123595506, -81.9101123595506,
  -80.8988764044944, -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944, 
    -80.8988764044944, -80.8988764044944, -80.8988764044944,
  -79.8876404494382, -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382, 
    -79.8876404494382, -79.8876404494382, -79.8876404494382,
  -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382, -78.876404494382, -78.876404494382, -78.876404494382, 
    -78.876404494382,
  -77.8651685393259, -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259, 
    -77.8651685393259, -77.8651685393259, -77.8651685393259,
  -76.8539325842697, -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697, 
    -76.8539325842697, -76.8539325842697, -76.8539325842697,
  -75.8426966292135, -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135, 
    -75.8426966292135, -75.8426966292135, -75.8426966292135,
  -74.8314606741573, -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573, 
    -74.8314606741573, -74.8314606741573, -74.8314606741573,
  -73.8202247191011, -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011, 
    -73.8202247191011, -73.8202247191011, -73.8202247191011,
  -72.8089887640449, -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449, 
    -72.8089887640449, -72.8089887640449, -72.8089887640449,
  -71.7977528089888, -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888, 
    -71.7977528089888, -71.7977528089888, -71.7977528089888,
  -70.7865168539326, -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326, 
    -70.7865168539326, -70.7865168539326, -70.7865168539326,
  -69.7752808988764, -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764, 
    -69.7752808988764, -69.7752808988764, -69.7752808988764,
  -68.7640449438202, -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202, 
    -68.7640449438202, -68.7640449438202, -68.7640449438202,
  -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764, -67.752808988764, -67.752808988764, -67.752808988764, 
    -67.752808988764,
  -66.7415730337079, -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079, 
    -66.7415730337079, -66.7415730337079, -66.7415730337079,
  -65.7303370786517, -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517, 
    -65.7303370786517, -65.7303370786517, -65.7303370786517,
  -64.7191011235955, -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955, 
    -64.7191011235955, -64.7191011235955, -64.7191011235955,
  -63.7078651685393, -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393, 
    -63.7078651685393, -63.7078651685393, -63.7078651685393,
  -62.6966292134831, -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831, 
    -62.6966292134831, -62.6966292134831, -62.6966292134831,
  -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427, -61.685393258427, -61.685393258427, -61.685393258427, 
    -61.685393258427,
  -60.6741573033708, -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708, 
    -60.6741573033708, -60.6741573033708, -60.6741573033708,
  -59.6629213483146, -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146, 
    -59.6629213483146, -59.6629213483146, -59.6629213483146,
  -58.6516853932584, -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584, 
    -58.6516853932584, -58.6516853932584, -58.6516853932584,
  -57.6404494382022, -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022, 
    -57.6404494382022, -57.6404494382022, -57.6404494382022,
  -56.6292134831461, -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461, 
    -56.6292134831461, -56.6292134831461, -56.6292134831461,
  -55.6179775280899, -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899, 
    -55.6179775280899, -55.6179775280899, -55.6179775280899,
  -54.6067415730337, -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337, 
    -54.6067415730337, -54.6067415730337, -54.6067415730337,
  -53.5955056179775, -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775, 
    -53.5955056179775, -53.5955056179775, -53.5955056179775,
  -52.5842696629214, -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214, 
    -52.5842696629214, -52.5842696629214, -52.5842696629214,
  -51.5730337078652, -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652, 
    -51.5730337078652, -51.5730337078652, -51.5730337078652,
  -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809, -50.561797752809, -50.561797752809, -50.561797752809, 
    -50.561797752809,
  -49.5505617977528, -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528, 
    -49.5505617977528, -49.5505617977528, -49.5505617977528,
  -48.5393258426966, -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966, 
    -48.5393258426966, -48.5393258426966, -48.5393258426966,
  -47.5280898876404, -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404, 
    -47.5280898876404, -47.5280898876404, -47.5280898876404,
  -46.5168539325843, -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843, 
    -46.5168539325843, -46.5168539325843, -46.5168539325843,
  -45.5056179775281, -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281, 
    -45.5056179775281, -45.5056179775281, -45.5056179775281,
  -44.4943820224719, -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719, 
    -44.4943820224719, -44.4943820224719, -44.4943820224719,
  -43.4831460674157, -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157, 
    -43.4831460674157, -43.4831460674157, -43.4831460674157,
  -42.4719101123596, -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596, 
    -42.4719101123596, -42.4719101123596, -42.4719101123596,
  -41.4606741573034, -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034, 
    -41.4606741573034, -41.4606741573034, -41.4606741573034,
  -40.4494382022472, -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472, 
    -40.4494382022472, -40.4494382022472, -40.4494382022472,
  -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191, -39.438202247191, -39.438202247191, -39.438202247191, 
    -39.438202247191,
  -38.4269662921348, -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348, 
    -38.4269662921348, -38.4269662921348, -38.4269662921348,
  -37.4157303370786, -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786, 
    -37.4157303370786, -37.4157303370786, -37.4157303370786,
  -36.4044943820225, -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225, 
    -36.4044943820225, -36.4044943820225, -36.4044943820225,
  -35.3932584269663, -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663, 
    -35.3932584269663, -35.3932584269663, -35.3932584269663,
  -34.3820224719101, -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101, 
    -34.3820224719101, -34.3820224719101, -34.3820224719101,
  -33.3707865168539, -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539, 
    -33.3707865168539, -33.3707865168539, -33.3707865168539,
  -32.3595505617978, -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978, 
    -32.3595505617978, -32.3595505617978, -32.3595505617978,
  -31.3483146067416, -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416, 
    -31.3483146067416, -31.3483146067416, -31.3483146067416,
  -30.3370786516854, -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854, 
    -30.3370786516854, -30.3370786516854, -30.3370786516854,
  -29.3258426966292, -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292, 
    -29.3258426966292, -29.3258426966292, -29.3258426966292,
  -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573, -28.314606741573, -28.314606741573, -28.314606741573, 
    -28.314606741573,
  -27.3033707865169, -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169, 
    -27.3033707865169, -27.3033707865169, -27.3033707865169,
  -26.2921348314607, -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607, 
    -26.2921348314607, -26.2921348314607, -26.2921348314607,
  -25.2808988764045, -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045, 
    -25.2808988764045, -25.2808988764045, -25.2808988764045,
  -24.2696629213483, -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483, 
    -24.2696629213483, -24.2696629213483, -24.2696629213483,
  -23.2584269662921, -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921, 
    -23.2584269662921, -23.2584269662921, -23.2584269662921,
  -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236, -22.247191011236, -22.247191011236, -22.247191011236, 
    -22.247191011236,
  -21.2359550561798, -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798, 
    -21.2359550561798, -21.2359550561798, -21.2359550561798,
  -20.2247191011236, -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236, 
    -20.2247191011236, -20.2247191011236, -20.2247191011236,
  -19.2134831460674, -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674, 
    -19.2134831460674, -19.2134831460674, -19.2134831460674,
  -18.2022471910112, -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112, 
    -18.2022471910112, -18.2022471910112, -18.2022471910112,
  -17.1910112359551, -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551, 
    -17.1910112359551, -17.1910112359551, -17.1910112359551,
  -16.1797752808989, -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989, 
    -16.1797752808989, -16.1797752808989, -16.1797752808989,
  -15.1685393258427, -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427, 
    -15.1685393258427, -15.1685393258427, -15.1685393258427,
  -14.1573033707865, -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865, 
    -14.1573033707865, -14.1573033707865, -14.1573033707865,
  -13.1460674157303, -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303, 
    -13.1460674157303, -13.1460674157303, -13.1460674157303,
  -12.1348314606742, -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742, 
    -12.1348314606742, -12.1348314606742, -12.1348314606742,
  -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618, -11.123595505618, -11.123595505618, -11.123595505618, 
    -11.123595505618,
  -10.1123595505618, -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618, 
    -10.1123595505618, -10.1123595505618, -10.1123595505618,
  -9.10112359550561, -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561, 
    -9.10112359550561, -9.10112359550561, -9.10112359550561,
  -8.08988764044943, -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943, 
    -8.08988764044943, -8.08988764044943, -8.08988764044943,
  -7.07865168539325, -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325, 
    -7.07865168539325, -7.07865168539325, -7.07865168539325,
  -6.06741573033707, -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707, 
    -6.06741573033707, -6.06741573033707, -6.06741573033707,
  -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809, -5.0561797752809, -5.0561797752809, -5.0561797752809, 
    -5.0561797752809,
  -4.04494382022472, -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472, 
    -4.04494382022472, -4.04494382022472, -4.04494382022472,
  -3.03370786516854, -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854, 
    -3.03370786516854, -3.03370786516854, -3.03370786516854,
  -2.02247191011236, -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236, 
    -2.02247191011236, -2.02247191011236, -2.02247191011236,
  -1.01123595505618, -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618, 
    -1.01123595505618, -1.01123595505618, -1.01123595505618,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618, 1.01123595505618, 1.01123595505618, 1.01123595505618, 
    1.01123595505618,
  2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236, 2.02247191011236, 2.02247191011236, 2.02247191011236, 
    2.02247191011236,
  3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854, 3.03370786516854, 3.03370786516854, 3.03370786516854, 
    3.03370786516854,
  4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472, 4.04494382022472, 4.04494382022472, 4.04494382022472, 
    4.04494382022472,
  5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809, 5.0561797752809, 5.0561797752809, 5.0561797752809, 
    5.0561797752809,
  6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707, 6.06741573033707, 6.06741573033707, 6.06741573033707, 
    6.06741573033707,
  7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325, 7.07865168539325, 7.07865168539325, 7.07865168539325, 
    7.07865168539325,
  8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943, 8.08988764044943, 8.08988764044943, 8.08988764044943, 
    8.08988764044943,
  9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561, 9.10112359550561, 9.10112359550561, 9.10112359550561, 
    9.10112359550561,
  10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618, 10.1123595505618, 10.1123595505618, 10.1123595505618, 
    10.1123595505618,
  11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618, 11.123595505618, 11.123595505618, 11.123595505618, 
    11.123595505618,
  12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742, 12.1348314606742, 12.1348314606742, 12.1348314606742, 
    12.1348314606742,
  13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303, 13.1460674157303, 13.1460674157303, 13.1460674157303, 
    13.1460674157303,
  14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865, 14.1573033707865, 14.1573033707865, 14.1573033707865, 
    14.1573033707865,
  15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427, 15.1685393258427, 15.1685393258427, 15.1685393258427, 
    15.1685393258427,
  16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989, 16.1797752808989, 16.1797752808989, 16.1797752808989, 
    16.1797752808989,
  17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551, 17.1910112359551, 17.1910112359551, 17.1910112359551, 
    17.1910112359551,
  18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112, 18.2022471910112, 18.2022471910112, 18.2022471910112, 
    18.2022471910112,
  19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674, 19.2134831460674, 19.2134831460674, 19.2134831460674, 
    19.2134831460674,
  20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236, 20.2247191011236, 20.2247191011236, 20.2247191011236, 
    20.2247191011236,
  21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798, 21.2359550561798, 21.2359550561798, 21.2359550561798, 
    21.2359550561798,
  22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236, 22.247191011236, 22.247191011236, 22.247191011236, 
    22.247191011236,
  23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921, 23.2584269662921, 23.2584269662921, 23.2584269662921, 
    23.2584269662921,
  24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483, 24.2696629213483, 24.2696629213483, 24.2696629213483, 
    24.2696629213483,
  25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045, 25.2808988764045, 25.2808988764045, 25.2808988764045, 
    25.2808988764045,
  26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607, 26.2921348314607, 26.2921348314607, 26.2921348314607, 
    26.2921348314607,
  27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169, 27.3033707865169, 27.3033707865169, 27.3033707865169, 
    27.3033707865169,
  28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573, 28.314606741573, 28.314606741573, 28.314606741573, 
    28.314606741573,
  29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292, 29.3258426966292, 29.3258426966292, 29.3258426966292, 
    29.3258426966292,
  30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854, 30.3370786516854, 30.3370786516854, 30.3370786516854, 
    30.3370786516854,
  31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416, 31.3483146067416, 31.3483146067416, 31.3483146067416, 
    31.3483146067416,
  32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977, 32.3595505617977, 32.3595505617977, 32.3595505617977, 
    32.3595505617977,
  33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539, 33.3707865168539, 33.3707865168539, 33.3707865168539, 
    33.3707865168539,
  34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101, 34.3820224719101, 34.3820224719101, 34.3820224719101, 
    34.3820224719101,
  35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663, 35.3932584269663, 35.3932584269663, 35.3932584269663, 
    35.3932584269663,
  36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225, 36.4044943820225, 36.4044943820225, 36.4044943820225, 
    36.4044943820225,
  37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787, 37.4157303370787, 37.4157303370787, 37.4157303370787, 
    37.4157303370787,
  38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348, 38.4269662921348, 38.4269662921348, 38.4269662921348, 
    38.4269662921348,
  39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191, 39.438202247191, 39.438202247191, 39.438202247191, 
    39.438202247191,
  40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472, 40.4494382022472, 40.4494382022472, 40.4494382022472, 
    40.4494382022472,
  41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034, 41.4606741573034, 41.4606741573034, 41.4606741573034, 
    41.4606741573034,
  42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596, 42.4719101123596, 42.4719101123596, 42.4719101123596, 
    42.4719101123596,
  43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157, 43.4831460674157, 43.4831460674157, 43.4831460674157, 
    43.4831460674157,
  44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719, 44.4943820224719, 44.4943820224719, 44.4943820224719, 
    44.4943820224719,
  45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281, 45.5056179775281, 45.5056179775281, 45.5056179775281, 
    45.5056179775281,
  46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843, 46.5168539325843, 46.5168539325843, 46.5168539325843, 
    46.5168539325843,
  47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404, 47.5280898876404, 47.5280898876404, 47.5280898876404, 
    47.5280898876404,
  48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966, 48.5393258426966, 48.5393258426966, 48.5393258426966, 
    48.5393258426966,
  49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528, 49.5505617977528, 49.5505617977528, 49.5505617977528, 
    49.5505617977528,
  50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809, 50.561797752809, 50.561797752809, 50.561797752809, 
    50.561797752809,
  51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652, 51.5730337078652, 51.5730337078652, 51.5730337078652, 
    51.5730337078652,
  52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213, 52.5842696629213, 52.5842696629213, 52.5842696629213, 
    52.5842696629213,
  53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775, 53.5955056179775, 53.5955056179775, 53.5955056179775, 
    53.5955056179775,
  54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337, 54.6067415730337, 54.6067415730337, 54.6067415730337, 
    54.6067415730337,
  55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899, 55.6179775280899, 55.6179775280899, 55.6179775280899, 
    55.6179775280899,
  56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461, 56.6292134831461, 56.6292134831461, 56.6292134831461, 
    56.6292134831461,
  57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022, 57.6404494382022, 57.6404494382022, 57.6404494382022, 
    57.6404494382022,
  58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584, 58.6516853932584, 58.6516853932584, 58.6516853932584, 
    58.6516853932584,
  59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146, 59.6629213483146, 59.6629213483146, 59.6629213483146, 
    59.6629213483146,
  60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708, 60.6741573033708, 60.6741573033708, 60.6741573033708, 
    60.6741573033708,
  61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427, 61.685393258427, 61.685393258427, 61.685393258427, 
    61.685393258427,
  62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831, 62.6966292134831, 62.6966292134831, 62.6966292134831, 
    62.6966292134831,
  63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393, 63.7078651685393, 63.7078651685393, 63.7078651685393, 
    63.7078651685393,
  64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955, 64.7191011235955, 64.7191011235955, 64.7191011235955, 
    64.7191011235955,
  65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517, 65.7303370786517, 65.7303370786517, 65.7303370786517, 
    65.7303370786517,
  66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079, 66.7415730337079, 66.7415730337079, 66.7415730337079, 
    66.7415730337079,
  67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764, 67.752808988764, 67.752808988764, 67.752808988764, 
    67.752808988764,
  68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202, 68.7640449438202, 68.7640449438202, 68.7640449438202, 
    68.7640449438202,
  69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764, 69.7752808988764, 69.7752808988764, 69.7752808988764, 
    69.7752808988764,
  70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326, 70.7865168539326, 70.7865168539326, 70.7865168539326, 
    70.7865168539326,
  71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888, 71.7977528089888, 71.7977528089888, 71.7977528089888, 
    71.7977528089888,
  72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045, 72.808988764045, 72.808988764045, 72.808988764045, 
    72.808988764045,
  73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011, 73.8202247191011, 73.8202247191011, 73.8202247191011, 
    73.8202247191011,
  74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573, 74.8314606741573, 74.8314606741573, 74.8314606741573, 
    74.8314606741573,
  75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135, 75.8426966292135, 75.8426966292135, 75.8426966292135, 
    75.8426966292135,
  76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697, 76.8539325842697, 76.8539325842697, 76.8539325842697, 
    76.8539325842697,
  77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259, 77.8651685393259, 77.8651685393259, 77.8651685393259, 
    77.8651685393259,
  78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382, 78.876404494382, 78.876404494382, 78.876404494382, 
    78.876404494382,
  79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382, 79.8876404494382, 79.8876404494382, 79.8876404494382, 
    79.8876404494382,
  80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944, 80.8988764044944, 80.8988764044944, 80.8988764044944, 
    80.8988764044944,
  81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506, 81.9101123595506, 81.9101123595506, 81.9101123595506, 
    81.9101123595506,
  82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067, 82.9213483146067, 82.9213483146067, 82.9213483146067, 
    82.9213483146067,
  83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629, 83.9325842696629, 83.9325842696629, 83.9325842696629, 
    83.9325842696629,
  84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191, 84.9438202247191, 84.9438202247191, 84.9438202247191, 
    84.9438202247191,
  85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753, 85.9550561797753, 85.9550561797753, 85.9550561797753, 
    85.9550561797753,
  86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315, 86.9662921348315, 86.9662921348315, 86.9662921348315, 
    86.9662921348315,
  87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876, 87.9775280898876, 87.9775280898876, 87.9775280898876, 
    87.9775280898876,
  88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438, 88.9887640449438, 88.9887640449438, 88.9887640449438, 
    88.9887640449438,
  89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719, 89.4943820224719, 89.4943820224719, 89.4943820224719, 
    89.4943820224719,
  90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 
    90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90 ;

 dx =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 dy =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 angle_dx =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 area =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;
}
