netcdf topog {
dimensions:
	nx = 360 ;
	ny = 200 ;
variables:
	double depth(ny, nx) ;
		depth:standard_name = "topographic depth at T-cell centers" ;
		depth:units = "meters" ;
data:

 depth =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 70, 253.361404418945, 
    253.361404418945, 253.361404418945, 305.484527587891, 341.096984863281, 
    625.089172363281, 702.910766601562, 683.282409667969, 666.132934570312, 
    566.239562988281, 456.478973388672, 456.478973388672, 448.196472167969, 
    455, 455, 455, 641.025512695312, 649.506164550781, 566.529724121094, 
    564.372741699219, 529.277099609375, 525, 525, 525, 452.484680175781, 
    458.936157226562, 458.936157226562, 451.466033935547, 471.123962402344, 
    439.039520263672, 462.933898925781, 480.040649414062, 557.98974609375, 
    566.638488769531, 566.638488769531, 502.514495849609, 395.754150390625, 
    395.754150390625, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    90, 140, 190, 230, 278.927978515625, 313.071350097656, 349.386352539062, 
    389.799438476562, 469.588500976562, 540.061584472656, 710.108276367188, 
    836.558532714844, 836.558532714844, 513.387145996094, 240.561416625977, 
    70, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 393.779937744141, 
    671.374389648438, 645.381042480469, 555, 555, 555, 625.089172363281, 
    764.700805664062, 729.532409667969, 666.132934570312, 566.239562988281, 
    456.478973388672, 461.591064453125, 448.196472167969, 455, 455, 455, 
    581.957702636719, 589.593017578125, 566.529724121094, 564.372741699219, 
    529.277099609375, 525, 525, 525, 452.484680175781, 458.936157226562, 
    466.627593994141, 451.466033935547, 441.517333984375, 425.785466617812, 
    453.429718017578, 480.040649414062, 566.638488769531, 566.638488769531, 
    752.81494140625, 735.182312011719, 811.403015136719, 922.524108886719, 
    1090.29431152344, 1090.29431152344, 1037.87707519531, 950.712585449219, 
    655.329162597656, 377.868743896484, 315, 120, 0, 0, 0, 0, 0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 200, 200, 200, 
    200, 200, 276.838012695312, 270.610395222517, 253.361404418945, 
    253.361404418945, 278.927978515625, 313.071350097656, 349.386352539062, 
    389.799438476562, 469.588500976562, 540.061584472656, 710.108276367188, 
    836.558532714844, 911.703369140625, 545.548278808594, 560.739196777344, 
    570.638916015625, 570.638916015625, 405.115844726562, 270.610395222517, 
    120, 110, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 393.779937744141, 
    645.381042480469, 645.381042480469, 555, 555, 555, 475, 502.862945556641, 
    502.862945556641, 476.903869628906, 400.195556640625, 316.587585449219, 
    372.031219482422, 401.529541015625, 455, 455, 455, 500.834838867188, 
    553.348571777344, 566.489196777344, 581.296997070312, 660.633178710938, 
    825.365234375, 1180.95568847656, 1478.68884277344, 1704.10205078125, 
    1878.22119140625, 1878.22119140625, 1732.318359375, 2087.44213867188, 
    2263.05078125, 2691.720703125, 2916.71533203125, 3078.25732421875, 
    3363.89404296875, 3356.07788085938, 3350.28540039062, 3466.79248046875, 
    3606.90063476562, 3624.53295898438, 3455.03051757812, 3552.80444335938, 
    3613.0478515625, 3574.12329101562, 3285.10668945312, 3256.55102539062, 
    2651.15991210938, 2386.88159179688, 1321.18334960938, 755.7919921875, 
    230, 140, 130, 110, 100, 90, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 
    200, 200, 200, 315, 543.88671875, 514.810119628906, 478.287963867188, 
    467.015777587891, 450.200378417969, 425.785466617812, 378.802062988281, 
    360, 294.462890625, 273.529113769531, 275.583374023438, 296.491394042969, 
    303.662811279297, 370.330291748047, 407.376525878906, 462.091278076172, 
    507.127319335938, 545.548278808594, 560.739196777344, 614.823791503906, 
    660.032897949219, 632.740783691406, 559.2138671875, 396.953247070312, 
    399.771759033203, 326.990295410156, 376.237579345703, 405.100372314453, 
    0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 90, 349.127227783203, 
    484.687072753906, 484.687072753906, 398.35986328125, 425.785466617812, 
    458.335906982422, 425.785466617812, 455, 455, 425.785466617812, 
    461.727447509766, 381.351470947266, 385.774627685547, 341.950958251953, 
    301.822479248047, 326.990295410156, 406.502563476562, 683.282409667969, 
    1252.83215332031, 1910.83435058594, 2191.85384798669, 2417.91015625, 
    2525.85034179688, 2733.93286132812, 3029.21850585938, 3041.10327148438, 
    3138.08959960938, 3171.37280273438, 3245.20043945312, 3540.50415039062, 
    3508.900390625, 3583.40698242188, 3640.20629882812, 3702.18188476562, 
    3651.04370117188, 3606.70092773438, 3725.0673828125, 3762.77319335938, 
    3795.36376953125, 3801.13525390625, 3869.6005859375, 3864.7890625, 
    3849.39428710938, 3844.142578125, 3924.37841796875, 3839.80859375, 
    3817.07177734375, 3725.72900390625, 3622.49975585938, 3475.25756835938, 
    2791.1845703125, 1870.03344726562, 1200.91442871094, 1192.88793945312, 
    819.087707519531, 473.113433837891, 441.202117919922, 388.126373291016, 
    388.126373291016, 230, 230, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 0, 0, 0, 200, 200, 315, 477.043304443359, 
    477.043304443359, 453.219696044922, 544.189208984375, 551.124328613281, 
    478.287963867188, 467.015777587891, 450.200378417969, 425.785466617812, 
    378.802062988281, 480.637054443359, 474.097717285156, 426.669372558594, 
    370.154968261719, 371.537628173828, 352.625915527344, 447.441925048828, 
    528.587646484375, 558.947021484375, 744.084777832031, 787.906860351562, 
    665.523498535156, 651.162109375, 667.357971191406, 667.357971191406, 
    747.587280273438, 923.585998535156, 923.585998535156, 611.835510253906, 
    604.615112304688, 562.673461914062, 562.673461914062, 522.4423828125, 
    347.727630615234, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 90, 140, 
    425.785466617812, 442.466430664062, 466.756195068359, 455, 455, 455, 455, 
    455, 429.319061279297, 425.785466617812, 386.934326171875, 
    390.988891601562, 449.432739257812, 788.671997070312, 1252.83215332031, 
    1910.83435058594, 2484.97119140625, 2893.2529296875, 2893.2529296875, 
    3135.48559570312, 3776.58056640625, 3886.513671875, 3918.4892578125, 
    3887.60766601562, 4005.93969726562, 4005.93969726562, 3986.43286132812, 
    3815.17944335938, 3779.66918945312, 3842.79541015625, 3998.97534179688, 
    3925.61743164062, 3908.76220703125, 4123.013671875, 4147.255859375, 
    4011.6728515625, 4096.5556640625, 4097.18896484375, 4038.5693359375, 
    4190.92919921875, 4177.61279296875, 4149.71826171875, 4124.390625, 
    4043.73608398438, 4027.92431640625, 3946.1533203125, 3925.6484375, 
    3921.86450195312, 3917.06127929688, 3847.74487304688, 3706.85131835938, 
    3706.85131835938, 3534.00732421875, 3161.671875, 2898.4033203125, 
    2931.53515625, 2976.1669921875, 2976.1669921875, 1953.28332519531, 
    1293.31567382812, 942.839303029559, 752.166198730469, 692.789672851562, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    470.156433105469, 470.156433105469, 130, 60, 60, 0, 0, 0, 0, -0, -0, -0, 
    -0, 0, -0, -0, 0, 0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 200, 360, 
    475.584625244141, 506.699859619141, 499.192993164062, 477.043304443359, 
    453.219696044922, 433.042846679688, 402.433135986328, 358.164398193359, 
    348.121124267578, 273.64208984375, 253.361404418945, 376.363647460938, 
    433.590576171875, 672.634765625, 836.252624511719, 977.149597167969, 
    1366.57861328125, 1787.79040527344, 2145.51684570312, 2335.1064453125, 
    2613.50805664062, 2828.27465820312, 2795.32299804688, 2765.18774414062, 
    2758.41088867188, 2743.02563476562, 2794.44653320312, 3065.78548661781, 
    3298.82299804688, 2923.783203125, 2448.35278320312, 2178.1806640625, 
    2178.1806640625, 2116.34765625, 1219.58276367188, 1010.98388671875, 
    594.427917480469, 328.744354248047, 120, 0, 0, 0, 0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    253.361404418945, 388.434295654297, 446.383087158203, 456.505737304688, 
    535.576843261719, 683.282409667969, 1019.00915527344, 1882.11401367188, 
    1819.87329101562, 1819.87329101562, 1286.38488769531, 604.795654296875, 
    587.180419921875, 683.282409667969, 1178.58068847656, 2484.97119140625, 
    3354.62280273438, 3688.7470703125, 3783.4970703125, 3787.27416992188, 
    3929.28149414062, 4004.40991210938, 4095.18334960938, 4219.64697265625, 
    4212.46728515625, 4197.943359375, 4198.46142578125, 4207.9814453125, 
    4215.0869140625, 4221.55712890625, 4212.76416015625, 4221.8701171875, 
    4237.58837890625, 4201.4423828125, 4182.82373046875, 4163.90185546875, 
    4189.22998046875, 4038.5693359375, 4144.91015625, 4152.17724609375, 
    4121.33642578125, 4212.880859375, 4210.19873046875, 4201.07666015625, 
    4175.69873046875, 4145.4697265625, 4075.30786132812, 4089.79150390625, 
    4100.673828125, 4125.56640625, 4069.76000976562, 3928.32495117188, 
    3865.92138671875, 3774.46606445312, 3632.576171875, 3655.435546875, 
    3341.38623046875, 3267.5087890625, 3201.10620117188, 3038.31005859375, 
    2758.41088867188, 2590.81884765625, 2387.99243164062, 2090.43823242188, 
    2142.17602539062, 2343.19848632812, 2241.88452148438, 1971.287109375, 
    1764.23596191406, 1454.45654296875, 1055.20068359375, 942.839303029559, 
    911.72265625, 889.461853027344, 863.093811035156, 850.199584960938, 
    789.079772949219, 842.674255371094, 852.9873046875, 863.308410644531, 
    880.477844238281, 904.889221191406, 898.118835449219, 913.220092773438, 
    756.595886230469, 506.711059570312, 381.929260253906, 40, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 281.439636230469, 338.740112304688, 
    338.740112304688, 294.462890625, 309.383575439453, 294.462890625, 
    312.565277099609, 331.474456787109, 380.938079833984, 370.497528076172, 
    302.059539794922, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, 
    0, 0, 200, 414.405670166016, 532.455444335938, 592.129211425781, 
    702.058166503906, 828.69384765625, 943.673400878906, 974.942504882812, 
    717.799865722656, 294.462890625, 255.369110107422, 90, 308.070892333984, 
    692.410217285156, 1240.05578613281, 1731.40795898438, 1974.732421875, 
    2368.20629882812, 2466.66776221529, 2907.00903320312, 3705.4931640625, 
    3705.4931640625, 3505.51025390625, 3533.82397460938, 3538.85668945312, 
    3462.86401367188, 3434.623046875, 3390.654296875, 3452.310546875, 
    3721.27612304688, 3931.17529296875, 3685.89599609375, 3555.61303710938, 
    3570.052734375, 3391.865234375, 3837.49877929688, 3939.57641601562, 
    3894.69921875, 3617.57861328125, 2868.96728515625, 2940.75903320312, 
    2166.62084960938, 401.556243896484, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    661.576293945312, 1847.98754882812, 2028.01293945312, 2177.63452148438, 
    2162.73583984375, 1835.923828125, 1715.58312988281, 1819.87329101562, 
    1819.87329101562, 1283.28967285156, 1213.70617675781, 1352.42797851562, 
    2031.31872558594, 2702.74145507812, 2896.41015625, 3671.12646484375, 
    3754.83520507812, 4035.37084960938, 4035.37084960938, 3952.63208007812, 
    4033.70678710938, 4164.36669921875, 4325.3994140625, 4314.982421875, 
    4235.94921875, 4195.072265625, 4162.583984375, 4256.767578125, 
    4275.32421875, 4298.716796875, 4287.9052734375, 4303.3759765625, 
    4317.94384765625, 4328.333984375, 4352.98486328125, 4314.47216796875, 
    4289.52587890625, 4265.13134765625, 4232.80908203125, 4183.5654296875, 
    4211.1171875, 4218.38330078125, 4231.5322265625, 4265.4091796875, 
    4234.43017578125, 4268.44775390625, 4285.521484375, 4281.31494140625, 
    4210.15380859375, 4229.607421875, 4179.3203125, 4174.134765625, 
    4225.2724609375, 4168.3896484375, 4078.7158203125, 4001.58178710938, 
    3790.982421875, 3663.25317382812, 3498.75317382812, 3353.36694335938, 
    3164.380859375, 3335.07397460938, 3374.45629882812, 3374.45629882812, 
    3304.5703125, 3088.55395507812, 2691.59643554688, 2691.59643554688, 
    2604.08520507812, 2347.18286132812, 1953.21069335938, 1747.7607421875, 
    1252.37072753906, 821.132873535156, 897.23095703125, 789.079772949219, 
    1017.75445556641, 1424.740234375, 1619.37915039062, 1647.68835449219, 
    1647.68835449219, 1647.68835449219, 1552.1513671875, 1254.10510253906, 
    899.144165039062, 921.160705566406, 921.160705566406, 442.385192871094, 
    451.422058105469, 451.422058105469, 170, 398.558288574219, 
    425.785466617812, 425.785466617812, 507.175354003906, 507.175354003906, 
    332.032318115234, 378.043762207031, 537.644287109375, 495.553629324057, 
    450.719116210938, 470.376647949219, 541.239990234375, 520.235229492188, 
    515.427062988281, 524.638977050781, 528.852844238281, 471.554534912109, 
    560, 560, 479.270538330078, 479.270538330078, 0, 0, 0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 253.361404418945, 414.405670166016, 
    580.953491210938, 774.6396484375, 737.9326171875, 1101.54602050781, 
    1530.7763671875, 1839.00744628906, 2112.47338867188, 2288.96606445312, 
    2267.34326171875, 2382.17529296875, 2560.90307617188, 2722.44555664062, 
    2904.08251953125, 3013.85717773438, 3250.82470703125, 3471.46630859375, 
    3804.03686523438, 3749.76733398438, 3814.62890625, 3897.30810546875, 
    3872.01391601562, 3872.6416015625, 3835.21899414062, 3881.75463867188, 
    3977.69555664062, 4109.66162109375, 4201.384765625, 4113.6552734375, 
    4023.04711914062, 4072.0087890625, 4124.634765625, 4022.5146484375, 
    4022.5146484375, 3993.4541015625, 4181.64111328125, 4250.787109375, 
    4331.42578125, 4331.6064453125, 4294.1396484375, 4038.94287109375, 
    3172.94921875, 2485.03955078125, 1886.56726074219, 771.988708496094, 
    278.569366455078, 278.569366455078, 0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, -0, 60, 60, 
    942.839303029559, 1682.87731933594, 2314.05395507812, 2314.05395507812, 
    2169.23876953125, 2113.47436523438, 2509.57421875, 2764.8408203125, 
    2822.65747070312, 3065.78548661781, 3117.54345703125, 3160, 3160, 3160, 
    3189.05322265625, 3869.78149414062, 3973.12646484375, 3973.12646484375, 
    4024.36108398438, 4047.10546875, 4047.10546875, 4035.37084960938, 
    4022.08471679688, 4033.70678710938, 4153.69482421875, 4197.00048828125, 
    4205.05908203125, 4273.4853515625, 4268.298828125, 4252.7978515625, 
    4254.33984375, 4240.9140625, 4356.71728515625, 4284.9423828125, 
    4272.45751953125, 4311.7412109375, 4383.93310546875, 4383.625, 
    4388.45751953125, 4359.28955078125, 4336.78076171875, 4309.52783203125, 
    4305, 4305, 4305, 4318.7294921875, 4321.60205078125, 4328.68310546875, 
    4290.36181640625, 4299.74755859375, 4302.9873046875, 4284.89990234375, 
    4329.00439453125, 4305.07275390625, 4356.91064453125, 4368.724609375, 
    4319.4169921875, 4207.24951171875, 4168.4921875, 4039.5712890625, 
    3938.60034179688, 3498.75317382812, 3353.36694335938, 3298.73388671875, 
    3335.07397460938, 3374.45629882812, 3374.45629882812, 3311.0693359375, 
    3160.61474609375, 2691.59643554688, 2691.59643554688, 2604.08520507812, 
    2680.22607421875, 2777.45654296875, 2933.0576171875, 3039.67944335938, 
    3292.64794921875, 3335.26977539062, 3335.26977539062, 3320.91552734375, 
    3221.20556640625, 3125.00122070312, 3291.39624023438, 3437.09912109375, 
    3588.47412109375, 3319.24438476562, 3181.84521484375, 3301.59399414062, 
    3301.59399414062, 3172.25512695312, 3264.74536132812, 3350.4375, 
    3350.4375, 3244.2275390625, 2597.63354492188, 1844.74035644531, 
    1236.87524414062, 916.291687011719, 1875.76171875, 2329.00830078125, 
    2406.9404296875, 2051.67749023438, 1468.45434570312, 1031.67529296875, 
    835.454284667969, 597.122863769531, 597.614074707031, 561.306945800781, 
    592.329284667969, 672.218994140625, 672.218994140625, 560, 560, 
    479.270538330078, 479.270538330078, 190, 0, 0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 0, 0, 370.154968261719, 551.57666015625, 
    580.953491210938, 738.946960449219, 1233.72204589844, 1975.87744140625, 
    2652.22216796875, 2825.05053710938, 2951.51611328125, 2927.82177734375, 
    3183.13500976562, 3312.97094726562, 3441.58154296875, 3543.30932617188, 
    3573.6376953125, 3567.68603515625, 3642.94775390625, 3756.50610351562, 
    3870.98364257812, 4068.689453125, 4192.92919921875, 4136.37890625, 
    4147.59423828125, 4165.1240234375, 4182.078125, 4171.779296875, 
    4237.0693359375, 4292.54052734375, 4306.005859375, 4403.5390625, 
    4461.22998046875, 4454.77734375, 4450.265625, 4433.830078125, 
    4358.6220703125, 4344.46630859375, 4399.50146484375, 4451.2080078125, 
    4444.9892578125, 4421.14501953125, 4455.212890625, 4532.17919921875, 
    4633.09912109375, 4607.9482421875, 4498.66357421875, 4032.37133789062, 
    2862.76928710938, 2244.88891601562, 1896.99938964844, 1446.50549316406, 
    731.054382324219, 520.916076660156, 495.553629324057, 485.388092041016, 
    294.462890625, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 190, 374.726104736328, 1068.52795410156, 
    1587.70288085938, 1761.97583007812, 1825.35913085938, 1983.79174804688, 
    2101.52978515625, 2358.80834960938, 2703.00732421875, 2702.76684570312, 
    2623.07958984375, 2169.23876953125, 2863.2197265625, 3188.7548828125, 
    3258.68530273438, 3360.85131835938, 3360.85131835938, 3360.85131835938, 
    3243.16430664062, 3161.19555664062, 3204.708984375, 3470.82446289062, 
    3869.78149414062, 4030.97680664062, 4044.48071289062, 4102.291015625, 
    4140.85888671875, 4047.10546875, 3957.70922851562, 4054.27880859375, 
    4026.486328125, 4026.486328125, 4189.3740234375, 4190.638671875, 
    4146.46142578125, 4026.81469726562, 4039.994140625, 4039.994140625, 
    4039.994140625, 4050, 4050, 4050, 4293.2373046875, 4248.90478515625, 
    4283.82470703125, 4359.28955078125, 4397.36083984375, 4397.36083984375, 
    4348.16796875, 4406.4892578125, 4379.23095703125, 4351.3818359375, 
    4330.828125, 4305, 4305, 4305, 4325.30810546875, 4341.1083984375, 
    4366.0048828125, 4384.275390625, 4395.9599609375, 4356.91064453125, 
    4374.05029296875, 4316.7197265625, 4338.71875, 4302.416015625, 
    4220.77099609375, 4017.71801757812, 3211.07446289062, 3648.41723632812, 
    3649.0498046875, 3521.05834960938, 3229.20263671875, 3229.20263671875, 
    2991.82250976562, 3559.03002929688, 3706.138671875, 3175.998046875, 
    2466.66776221529, 2903.63793945312, 2995.00927734375, 2995.00927734375, 
    3528.27807617188, 3721.27612304688, 3891.89721679688, 4010.443359375, 
    3612.61987304688, 3644.96142578125, 3750.9560546875, 3871.8974609375, 
    3912.39501953125, 3932.5810546875, 4035.083984375, 3877.099609375, 
    4031.7548828125, 4066.82861328125, 4212.3017578125, 4333.38330078125, 
    4229.166015625, 4214.41162109375, 4340.25146484375, 4319.873046875, 
    4332.662109375, 4362.02880859375, 3809.29174804688, 3840.912109375, 
    4005.3857421875, 4025.70849609375, 3227.58764648438, 3269.77685546875, 
    3269.77685546875, 2743.57958984375, 2466.66776221529, 2365.03735351562, 
    2536.638671875, 2466.66776221529, 1513.06506347656, 1029.31298828125, 
    845.613037109375, 636.124389648438, 620.577514648438, 391.155364990234, 
    190, 200, 200, 200, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 
    482.893127441406, 551.57666015625, 555.61328125, 646.677734375, 
    1329.76025390625, 2143.92846679688, 2652.22216796875, 2825.05053710938, 
    3028.27856445312, 3223.11767578125, 3516.03051757812, 3651.63989257812, 
    3507.36694335938, 3590.97412109375, 3916.91918945312, 3919.80932617188, 
    3912.24340820312, 3937.302734375, 3945.78051757812, 4091.71411132812, 
    4294.265625, 4276.88720703125, 4254.09619140625, 4271.24072265625, 
    4364.6640625, 4510.6923828125, 4419.18185522252, 4479.05029296875, 
    4542.0361328125, 4544.45068359375, 4595.2314453125, 4605.501953125, 
    4627.509765625, 4648.80615234375, 4607.4404296875, 4651.12939453125, 
    4643.826171875, 4680.572265625, 4656.943359375, 4638.48095703125, 
    4595.26708984375, 4632.8681640625, 4640.66748046875, 4702.84228515625, 
    4674.24169921875, 4757.76025390625, 4674.3349609375, 4527.6259765625, 
    4334.8056640625, 3612.70190429688, 2950.25854492188, 3003.30078125, 
    2952.767578125, 2796.38745117188, 1984.68054199219, 2714.95336914062, 
    2961.01953125, 3051.44677734375, 2654.78466796875, 2093.35327148438, 
    1590.93969726562, 2209.49291992188, 2325.01928710938, 2295.11279296875, 
    2330.29931640625, 1974.32141113281, 1601.46130371094, 1599.10827636719, 
    1817.56262207031, 1817.56262207031, 1240.76452636719, 310.411529541016, 
    220, 120, 150, 190, 425.785466617812, 639.720336914062, 1478.68884277344, 
    1956.08947753906, 1956.08947753906, 2129.50048828125, 2594.5205078125, 
    2929.12939453125, 2846.72680664062, 2520.291015625, 2037.18017578125, 
    1375.06274414062, 619.856750488281, 0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 
    0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 80, 80, 80, 80, 
    -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, -0, 
    0, 306.650299072266, 331.5927734375, 545.521301269531, 1103.45166015625, 
    1588.18908691406, 1942.33386230469, 2143.31079101562, 2352.16845703125, 
    2352.16845703125, 1761.97583007812, 1825.35913085938, 1983.79174804688, 
    2101.52978515625, 2358.80834960938, 2744.2890625, 2999.5751953125, 
    2961.00512695312, 2961.4951171875, 2961.4951171875, 3314.04248046875, 
    3481.8623046875, 3474.44848632812, 3360.85131835938, 3360.85131835938, 
    3243.16430664062, 3161.19555664062, 3142.09521484375, 3470.82446289062, 
    3686.3876953125, 3663.40502929688, 4046.50854492188, 4129.60595703125, 
    4155.24560546875, 3736.71215820312, 3901.70825195312, 3731.44555664062, 
    3755.33276367188, 3721.27612304688, 3874.41650390625, 4009.83447265625, 
    3786.72216796875, 3930.00048828125, 3806.18969726562, 3721.27612304688, 
    3835.958984375, 4050, 4050, 4050, 4067.96997070312, 4170.00439453125, 
    4239.703125, 4181.79638671875, 4397.36083984375, 4397.36083984375, 
    4348.16796875, 4379.23095703125, 4379.23095703125, 4373.40966796875, 
    4326.77392578125, 4305, 4305, 4305, 4303.619140625, 4335, 4335, 
    4362.0830078125, 4346.806640625, 4316.66259765625, 4326.52001953125, 
    4300.17919921875, 4343.755859375, 4348.18994140625, 4274.8544921875, 
    4215.7978515625, 4185.1953125, 4065.89147763595, 3855.546875, 
    3839.05151367188, 3989.52172851562, 4016.80053710938, 4065.89147763595, 
    4116.49609375, 4284.84765625, 4264.44921875, 4020.9599609375, 
    4054.04321289062, 4022.150390625, 4044.6220703125, 4099.830078125, 
    4262.958984375, 4268.97265625, 4249.2783203125, 4093.34033203125, 
    3983.974609375, 3945.0751953125, 4018.36987304688, 4234.92724609375, 
    4066.20166015625, 4317.21240234375, 4364.8759765625, 4276.27880859375, 
    4319.22998046875, 4328.50732421875, 4444.57080078125, 4490.37451171875, 
    4476.64208984375, 4521.31396484375, 4343.80419921875, 4463.87353515625, 
    4442.88623046875, 4419.18185522252, 4291.77197265625, 4374.53515625, 
    4065.89147763595, 3227.58764648438, 3876.8447265625, 3844.32861328125, 
    3721.27612304688, 3544.96411132812, 3575.71142578125, 3611.59106445312, 
    3611.59106445312, 3501.69799804688, 3600.78784179688, 3600.78784179688, 
    3522.41650390625, 3562.2607421875, 3343.58813476562, 2270.78100585938, 
    524.135009765625, 551.836181640625, 430.078308105469, 448.098388671875, 
    315.688293457031, 315.688293457031, 279.634033203125, -0, -0, -0, -0, 0, 
    0, 0, 0, 0, 482.893127441406, 539.531799316406, 495.553629324057, 
    463.441131591797, 1371.28747558594, 2085.34594726562, 2202.68994140625, 
    2807.71728515625, 3028.27856445312, 3223.11767578125, 3387.2978515625, 
    3418.95141601562, 3507.36694335938, 3590.97412109375, 3841.46655273438, 
    4027.68481445312, 4142.12158203125, 4260.79345703125, 4205.142578125, 
    4309.07958984375, 4335.13037109375, 4323.54931640625, 4435.54443359375, 
    4467.38427734375, 4472.310546875, 4442.689453125, 4444.10302734375, 
    4530.12353515625, 4587.23583984375, 4612.71240234375, 4632.0478515625, 
    4662.17578125, 4697.36572265625, 4722.55224609375, 4817.38525390625, 
    4820.83154296875, 4800.390625, 4789.46826171875, 4843.02734375, 
    4835.806640625, 4762.03076171875, 4791.63525390625, 4836.6259765625, 
    4757.76806640625, 4784.34423828125, 4810.46142578125, 4847.04150390625, 
    4887.00732421875, 4851.16064453125, 4540.43994140625, 4142.0654296875, 
    4026.30810546875, 3657.88525390625, 3408.85913085938, 3653.576171875, 
    3695.99633789062, 3900.02465820312, 4037.02880859375, 4029.56518554688, 
    4197.62353515625, 4241.4873046875, 4350.30859375, 4033.34912109375, 
    3628.71411132812, 3302.31103515625, 3328.40356445312, 3416.46948242188, 
    3503.77880859375, 3397.4765625, 3282.78540039062, 2815.24731445312, 
    1738.65734863281, 2163.03833007812, 2824.265625, 2983.01586914062, 
    3360.85571289062, 3360.85571289062, 3619.57495117188, 3619.57495117188, 
    3822.19018554688, 3762.21801757812, 3974.07592773438, 3816.94311523438, 
    3506.07055664062, 3494.10083007812, 3653.02685546875, 3584.99609375, 
    3655.80859375, 3270.66235351562, 2766.41943359375, 1801.34167480469, 
    335.664855957031, 240.762069702148, 0, 0, 220, 480, 755, 755, 
    326.990295410156, 326.990295410156, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 160, 444.9716796875, 568.222106933594, 568.222106933594, 
    451.431610107422, 410.269195556641, 341.01806640625, 295.040374755859, 
    -0, -0,
  357.184204101562, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 200, 
    315.078186035156, 581.105041503906, 738.803771972656, 715.2412109375, 
    610.024780273438, 627.470520019531, 525.640502929688, 525.640502929688, 
    462.864898681641, 1662.95068359375, 2435.50463867188, 2475.19018554688, 
    2543.57080078125, 2563.26171875, 2352.16845703125, 2386.69067382812, 
    991.139587402344, 1549.96508789062, 1658.74084472656, 1602.70922851562, 
    2073.37670898438, 2744.2890625, 2961.00512695312, 2961.00512695312, 
    3158.26293945312, 3187.62963867188, 3314.04248046875, 3542.62060546875, 
    3675.91015625, 3593.40649414062, 3621.79174804688, 3243.16430664062, 
    3150, 3142.09521484375, 3707.60595703125, 3663.40502929688, 
    3663.40502929688, 3680.20703125, 3273.12255859375, 3227.53393554688, 
    3201.21704101562, 3590.7890625, 3626.69799804688, 3419.42797851562, 
    3775.31762695312, 3786.3173828125, 3818.27783203125, 3840.77294921875, 
    3699.20874023438, 3513.81372070312, 3774.23071289062, 3962.87939453125, 
    3915.76977539062, 3972.38354492188, 3914.30004882812, 3952.650390625, 
    4055.24609375, 4055, 4055.72265625, 4255.86474609375, 4202.06201171875, 
    4253.39013671875, 4228.27685546875, 4159.1484375, 4173.89306640625, 
    4119.833984375, 4010, 4010, 4065.89147763595, 4125.15625, 
    4016.08251953125, 4287.56591796875, 4227.32666015625, 4316.66259765625, 
    4385.6904296875, 4335.337890625, 4426.30224609375, 4524.8115234375, 
    4420.17041015625, 4430.19482421875, 4452.17138671875, 4322.11865234375, 
    4306.931640625, 4357.794921875, 4362.80224609375, 4326.37744140625, 
    4254.01171875, 4184.2236328125, 4320.00146484375, 4287.73486328125, 
    4326.5556640625, 4387.521484375, 4386.513671875, 4388.85498046875, 
    4390.79833984375, 4452.890625, 4472.9638671875, 4490.9140625, 
    4407.49072265625, 4367.4677734375, 4276.28271484375, 4149.9521484375, 
    4089.17041015625, 4299.93359375, 4543.1376953125, 4606.69873046875, 
    4625.71923828125, 4700.2939453125, 4620.42041015625, 4625.55419921875, 
    4622.01708984375, 4630.03125, 4616.46728515625, 4605.22216796875, 
    4547.21875, 4548.26611328125, 4540.4921875, 4537.17041015625, 
    4539.3671875, 4468.20263671875, 4652.05517578125, 4280.5205078125, 
    4209.58203125, 4211.5478515625, 4241.18408203125, 4122.7119140625, 
    4180.7705078125, 4240.11083984375, 4175.298828125, 4176.34912109375, 
    4074.89501953125, 4093.775390625, 4107.25146484375, 3806.89184570312, 
    3474.84228515625, 3247.19384765625, 3251.38745117188, 2735.4677734375, 
    430.078308105469, 433.444030761719, 433.444030761719, 433.444030761719, 
    279.634033203125, -0, -0, -0, -0, -0, 0, 0, 0, 0, 392.230560302734, 
    509.845123291016, 534.733947753906, 588.047546386719, 1325.79724121094, 
    2085.34594726562, 2579.62524414062, 2975.775390625, 3134.197265625, 
    3317.11303710938, 3630.61376953125, 3709.59692382812, 3835.72021484375, 
    3869.45654296875, 3997.67919921875, 4047.7060546875, 4079.00854492188, 
    4177.744140625, 4310.16650390625, 4318.5986328125, 4371.45361328125, 
    4454.7998046875, 4474.84130859375, 4506.8447265625, 4614.8681640625, 
    4554.0068359375, 4570.2099609375, 4601.03466796875, 4594, 4597.75, 
    4658.8583984375, 4690.9873046875, 4733.0380859375, 4758.47119140625, 
    4842.97119140625, 4942.048828125, 4899.63525390625, 4867.71875, 
    4883.603515625, 4913.40673828125, 4876.1376953125, 4872.82666015625, 
    4960.16015625, 4974.974609375, 4911.6376953125, 4792.36962890625, 
    4915.3232421875, 4894.0703125, 4876.18359375, 4804.25048828125, 
    4727.29296875, 4915.9599609375, 4887.654296875, 4841.345703125, 
    4826.087890625, 4678.3134765625, 4454.552734375, 4306.34814453125, 
    4594.177734375, 4642.61279296875, 4241.4873046875, 4241.4873046875, 
    4033.34912109375, 3610.458984375, 4010.763671875, 4193.67041015625, 
    4228.21875, 4164.4365234375, 3902.42797851562, 3599.97265625, 
    2864.47314453125, 2468.6904296875, 3262.94677734375, 3325.61962890625, 
    3488.69213867188, 4070.18041992188, 4122.95361328125, 4382.85302734375, 
    4382.85302734375, 4220.01513671875, 4130.19287109375, 4387.09033203125, 
    4387.09033203125, 4324.697265625, 4227.94091796875, 4083.20458984375, 
    3971.0029296875, 3968.78051757812, 3874.49340820312, 3799.29760742188, 
    3562.439453125, 2860.31909179688, 1062.32312011719, 1130.1767578125, 
    2652.15161132812, 3374.93481445312, 3176.8408203125, 3410.83154296875, 
    3410.83154296875, 3226.15747070312, 2654.33056640625, 2654.33056640625, 
    1697.18078613281, 808.351013183594, 334.360778808594, 294.462890625, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 170, 
    326.990295410156, 326.990295410156, 326.990295410156, 253.361404418945, 
    270.610395222517, 307.885650634766, 547.565673828125, 568.222106933594, 
    568.222106933594, 451.431610107422, 410.269195556641, 341.01806640625, 
    295.040374755859, 310.406433105469, 428.268646240234,
  468.303649902344, 304.436859130859, 210, 150, 150, 0, -0, 0, 0, 220, 220, 
    140, 120, 60, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 
    -0, -0, -0, -0, -0, -0, 0, 391.194396972656, 473.844543457031, 
    473.844543457031, 385.810302734375, 120, 110, 130, 130, -0, -0, 80, 80, 
    80, -0, -0, -0, -0, -0, -0, -0, -0, 40, 277.445556640625, 294.462890625, 
    355.489166259766, 510.220550537109, 619.773193359375, 622.774841308594, 
    301.804107666016, 271.7666015625, 537.80224609375, 537.80224609375, 
    620.522338867188, 803.625015916513, 849.296447753906, 1284.23803710938, 
    1459.00268554688, 1459.00268554688, 2228.77978515625, 2618.36791992188, 
    2667.84790039062, 2851.34838867188, 2758.41088867188, 2643.0869140625, 
    2554.83984375, 830.093994140625, 2062.60083007812, 2468.2587890625, 
    2665.580078125, 2719.18505859375, 2876.54296875, 3045, 3045, 
    3001.93530273438, 3252.37866210938, 3168.18408203125, 3286.86596679688, 
    3223.70263671875, 3410.20849609375, 3593.40649414062, 3638.2431640625, 
    3510.8515625, 3065.78548661781, 2719.0419921875, 2719.0419921875, 
    2352.37548828125, 2801.53125, 2856.853515625, 3257.14428710938, 
    3166.67309570312, 3149.13452148438, 3088.39477539062, 3046.60400390625, 
    3261.73608398438, 3400.21118164062, 3630.68823242188, 3624.32495117188, 
    3624.4677734375, 3574.6513671875, 3574.6513671875, 3588.13452148438, 
    3721.27612304688, 3816.10375976562, 3915.76977539062, 3937.57470703125, 
    4027.58276367188, 3935.84912109375, 3961.17211914062, 4004.09155273438, 
    4055.72265625, 4206.47119140625, 4116.115234375, 4243.41748046875, 
    4256.9697265625, 4185, 4270.49462890625, 4210.5390625, 4010, 4010, 
    4011.36303710938, 4011.36303710938, 4016.08251953125, 4180.4189453125, 
    4271.24267578125, 4245.13623046875, 4236.61474609375, 4359.96728515625, 
    4578.28662109375, 4593.97900390625, 4616.95361328125, 4589.6318359375, 
    4653.93798828125, 4655.10986328125, 4601.703125, 4582.22900390625, 
    4642.462890625, 4562.4931640625, 4439.6044921875, 4458.56787109375, 
    4508.1416015625, 4551.74755859375, 4580.03759765625, 4667.97265625, 
    4717.56396484375, 4716.50830078125, 4718.12255859375, 4703.53515625, 
    4761.00927734375, 4793.8828125, 4828.98486328125, 4744.345703125, 
    4710.71533203125, 4541.5341796875, 4559.0810546875, 4588.7080078125, 
    4612.078125, 4704.4267578125, 4807.74609375, 4867.70458984375, 
    4814.30810546875, 4755.57568359375, 4753.154296875, 4738.7861328125, 
    4669.99169921875, 4695.142578125, 4744.9921875, 4723.91552734375, 
    4732.24951171875, 4672.00439453125, 4707.3564453125, 4737.0419921875, 
    4744.65380859375, 4280.5205078125, 4551.2744140625, 4486.96142578125, 
    4446.64892578125, 4438.1552734375, 4469.97509765625, 4493.181640625, 
    4433.97412109375, 4321.8291015625, 4255.00439453125, 4245.65625, 
    4106.09765625, 4007.94775390625, 3849.17456054688, 3510.30151367188, 
    3346.75537109375, 3490.90551757812, 3490.90551757812, 3362.21362304688, 
    1245.48034667969, 517.233947753906, 407.678558349609, 407.678558349609, 
    200, 40, -0, -0, 0, -0, 0, 0, 392.230560302734, 392.230560302734, 
    381.6904296875, 588.047546386719, 876.56689453125, 1745.64147949219, 
    2579.62524414062, 2975.775390625, 3134.197265625, 3317.11303710938, 
    3593.95385742188, 3917.7275390625, 3961.07055664062, 4140.5732421875, 
    4295.26708984375, 4285.7451171875, 4560, 4560, 4560, 4569.1748046875, 
    4568.587890625, 4738.677734375, 4589.9833984375, 4698.3505859375, 
    4646.17431640625, 4677.7861328125, 4691.6357421875, 4716.59716796875, 
    4731.7275390625, 4753.224609375, 4779.07571895829, 4816.7783203125, 
    4824.50537109375, 4838.01904296875, 4868.681640625, 4888.83837890625, 
    4902.7294921875, 4927.142578125, 4913.46826171875, 4949.23095703125, 
    4965.91455078125, 4976.90283203125, 5014.9736328125, 4987.29443359375, 
    4994.87451171875, 4998.7880859375, 5002.0908203125, 5004.74560546875, 
    4974.61376953125, 5062.47705078125, 5009.4658203125, 4945.4365234375, 
    4889.498046875, 4932.04931640625, 4861.11572265625, 4779.07571895829, 
    4601.28271484375, 4658.5791015625, 4717.98681640625, 4425, 
    3797.82885742188, 4046.53149414062, 3803.86401367188, 3667.23681640625, 
    4010.763671875, 4209.443359375, 4193.67041015625, 4283.2734375, 
    4270.734375, 3743.52294921875, 3548.97729492188, 3238.0693359375, 
    3287.21337890625, 3325.61962890625, 3680.501953125, 4154.181640625, 
    4349.8759765625, 4676.39013671875, 4684.87548828125, 4623.6494140625, 
    4599.3369140625, 4482.41552734375, 4604.40771484375, 4640.0283203125, 
    4594.7529296875, 4439.1162109375, 4419.18185522252, 4515.5302734375, 
    4296.53076171875, 4208.7275390625, 4187.3818359375, 3995.3388671875, 
    3373.0556640625, 1281.23913574219, 2696.9853515625, 4276.7080078125, 
    4419.18185522252, 4568.50732421875, 4527.04541015625, 4475.251953125, 
    4322.74658203125, 3815.58056640625, 3396.51025390625, 2947.05126953125, 
    2566.73779296875, 2466.66776221529, 1767.408203125, 1038.24133300781, 
    580.953491210938, 387.778839111328, -0, -0, -0, -0, -0, -0, -0, 
    432.559906005859, 702.638244628906, 1648.00842285156, 1676.32397460938, 
    1676.32397460938, 1708.75866699219, 2330.2568359375, 2437.85009765625, 
    2437.85009765625, 2111.76635742188, 2191.85384798669, 2191.85384798669, 
    1758.19494628906, 1758.19494628906, 1494.58935546875, 1284.02331542969, 
    1853.15869140625, 2373.84497070312, 2371.67016601562, 2298.98876953125, 
    2172.9609375, 1427.36608886719, 844.796020507812,
  2864.57495117188, 2163.88598632812, 2213.81103515625, 2359.0146484375, 
    2509.72802734375, 2703.48999023438, 2360.74145507812, 2238.72534179688, 
    2146.09057617188, 1963.53796386719, 1337.38012695312, 862.46484375, 
    510.071166992188, 425.785466617812, 299.707183837891, 0, -0, -0, 0, 0, 
    -0, 0, 0, 40, 240.561416625977, 327.056549072266, 669.441162109375, 
    669.441162109375, 560.386413574219, 580.953491210938, 803.625015916513, 
    920.105651855469, 920.105651855469, 541.93310546875, 541.93310546875, 
    440.315216064453, 374.443389892578, 709.050170898438, 709.050170898438, 
    1070.97009277344, 1601.43188476562, 1478.68884277344, 1193.41381835938, 
    1193.41381835938, 1156.58386230469, 560.070190429688, 387.852355957031, 
    387.852355957031, 383.570251464844, 258.796752929688, 619.186340332031, 
    619.186340332031, 542.29638671875, 542.29638671875, 294.462890625, 
    439.981353759766, 580.953491210938, 907.549438476562, 896.270690917969, 
    1186.69384765625, 1468.04846191406, 1586.48083496094, 1957.51220703125, 
    2327.28076171875, 2598.6416015625, 2636.55639648438, 2636.55639648438, 
    2982.78686523438, 2758.41088867188, 2679.64086914062, 2582.2880859375, 
    2523.51196289062, 2672.75317382812, 2672.75317382812, 3001.83227539062, 
    3001.83227539062, 2976.578125, 2904.17138671875, 2944.849609375, 
    2758.41088867188, 2699.02294921875, 2498.58422851562, 2874.892578125, 
    2862.04296875, 3051.29931640625, 3051.29931640625, 3051.244140625, 
    3021.07861328125, 3045, 3045, 3001.93530273438, 3231.61938476562, 
    3272.88623046875, 3243.95532226562, 3223.70263671875, 3364.04150390625, 
    3510, 3510, 3510, 2615, 2615, 2615, 2399.38330078125, 2493.11450195312, 
    2736.87744140625, 2516.49584960938, 2586.95385742188, 3025, 3025, 
    2939.43334960938, 2999.99267578125, 3004.61669921875, 3046.02392578125, 
    2980.42602539062, 3181.72607421875, 3438.4375, 3483.43872070312, 
    3588.13452148438, 3856.708984375, 3927.689453125, 3907.44702148438, 
    3937.57470703125, 3937.57470703125, 4048.81079101562, 3935.84912109375, 
    3835.44165039062, 3916.69799804688, 4005.80249023438, 3935.81274414062, 
    4100.4609375, 4195.52197265625, 4185, 4037.42602539062, 4054.66821289062, 
    3929.71313476562, 3983.61206054688, 4185, 4185, 4185, 4204.08642578125, 
    4164.9462890625, 4357.30419921875, 4249.9716796875, 4359.96728515625, 
    4583.67529296875, 4506.50830078125, 4659.00830078125, 4741.7314453125, 
    4779.07571895829, 4779.07571895829, 4711.30810546875, 4736.62353515625, 
    4699.35888671875, 4791.828125, 4779.61572265625, 4841.23095703125, 
    4793.6455078125, 4806.7900390625, 4829.52783203125, 4854.60791015625, 
    4892.6357421875, 4901.908203125, 4908.18115234375, 4878.2626953125, 
    4908.41162109375, 4867.4404296875, 4900.10546875, 4928.87451171875, 
    4919.44189453125, 4838.48828125, 4828.3154296875, 4789.923828125, 
    4819.08740234375, 4829.61474609375, 4967.109375, 4902.55126953125, 
    4907.72607421875, 4902.76171875, 4884.42626953125, 4880.18896484375, 
    4852.19873046875, 4815.34521484375, 4897.8525390625, 4818.89404296875, 
    4751.6611328125, 4752.8388671875, 4671.73291015625, 4671.73291015625, 
    4579.025390625, 4185, 4599.33203125, 4603.8486328125, 4548.9013671875, 
    4544.63330078125, 4509.556640625, 4501.09521484375, 4480.7255859375, 
    4336.20068359375, 4285.26220703125, 4202.56591796875, 4151.89111328125, 
    4041.95288085938, 4036.890625, 4043.34350585938, 4013.49438476562, 
    3632.89575195312, 3654.38671875, 3579.06005859375, 3307.32202148438, 
    3070.18408203125, 1385.59594726562, 425.785466617812, 200, 200, 60, 60, 
    -0, -0, 0, 0, 50, 370.154968261719, 381.6904296875, 384.316619873047, 
    451.619140625, 665.848449707031, 1796.32446289062, 2466.66776221529, 
    2931.57739257812, 3336.77319335938, 3711.17529296875, 3989.1259765625, 
    4036.1767578125, 4249.18505859375, 4301.0966796875, 4428.14404296875, 
    4528.1982421875, 4608.130859375, 4586.53466796875, 4642.5361328125, 
    4636.798828125, 4723.24755859375, 4745.84130859375, 4745.84130859375, 
    4762.4912109375, 4798.15869140625, 4806.39208984375, 4828.74462890625, 
    4842.232421875, 4877.06494140625, 4876.08349609375, 4890.65576171875, 
    4877.6357421875, 4913.23388671875, 4921.62451171875, 4970.49462890625, 
    4982.39892578125, 5053.623046875, 5052.7373046875, 4961.310546875, 
    4962.13037109375, 5006.921875, 5110.80615234375, 5082.68505859375, 
    5026.98583984375, 5111.73095703125, 5055.318359375, 5122.7041015625, 
    5117.333984375, 5055.3662109375, 5004.671875, 5019.4404296875, 
    4952.10986328125, 5000.22900390625, 5022.6142578125, 5020.8623046875, 
    4905.2431640625, 4891.43505859375, 4994.986328125, 4125.73876953125, 
    3205.376953125, 2943.3115234375, 2528.42797851562, 3123.5732421875, 
    3698.79370117188, 4244.87353515625, 4193.67041015625, 4239.85400390625, 
    4239.85400390625, 4377.6806640625, 4274.0224609375, 3909.1826171875, 
    3388.42333984375, 3367.28173828125, 3240.11694335938, 3513.79467773438, 
    3668.77026367188, 4614.53125, 4820.462890625, 4943.74169921875, 
    4860.3134765625, 4798.177734375, 4728.15380859375, 4795.216796875, 
    4884.06396484375, 4889.93701171875, 4829.64697265625, 4839.81982421875, 
    4793.68505859375, 4791.58544921875, 4785.09033203125, 4425.2705078125, 
    3566.54931640625, 3072.78637695312, 2696.9853515625, 4109.974609375, 
    4603.61181640625, 4779.07571895829, 4779.07571895829, 4737.98486328125, 
    4599.2509765625, 4352.6181640625, 3991.78466796875, 3628.42553710938, 
    3642.85717773438, 3479.8603515625, 3073.2412109375, 2532.13916015625, 
    2084.11181640625, 2346.6513671875, 2346.6513671875, 1764.47985839844, 
    1639.72045898438, 564.223999023438, 1051.26098632812, 2010.09924316406, 
    2332.03784179688, 2964.96411132812, 3426.97045898438, 3647.57666015625, 
    3741.11328125, 3887.6923828125, 3644.18310546875, 3467.49975585938, 
    2962.96142578125, 2801.84887695312, 3044.85278320312, 3044.85278320312, 
    2837.34594726562, 2662.82861328125, 2947.92260742188, 2965.24829101562, 
    2956.1259765625, 2993.83911132812, 2993.83911132812, 3257.45263671875, 
    3284.52221679688, 3284.52221679688, 3420.83178710938, 3391.91870117188,
  3647.92309570312, 3636.81591796875, 3475, 3475, 3556.7314453125, 
    3524.123046875, 3502.26879882812, 3368.27783203125, 3474.58862304688, 
    3526.8603515625, 3364.92431640625, 3054.83911132812, 2812.35791015625, 
    2492.17407226562, 1995.05810546875, 1006.36633300781, 742.55517578125, 
    413.826324462891, 413.826324462891, 391.662170410156, 90, 
    582.533081054688, 1422.44995117188, 1318.3603515625, 1961.06274414062, 
    1961.06274414062, 2603.166015625, 3114.99755859375, 3135.46166992188, 
    3112.201171875, 2832.56469726562, 2800.998046875, 2299.37963867188, 
    2302.15869140625, 1969.90783691406, 2059.48315429688, 2242.66577148438, 
    2580.33764648438, 2964.8486328125, 3083.36376953125, 3319.7919921875, 
    3154.35888671875, 3035.966796875, 2965.22485351562, 2973.90258789062, 
    3031.9404296875, 3031.9404296875, 2960.44970703125, 2521.09252929688, 
    2312.361328125, 1887.63903808594, 1887.63903808594, 1632.32995605469, 
    1869.41455078125, 2592.65771484375, 2643.27026367188, 2643.27026367188, 
    2998.162109375, 3206.18725585938, 3313.63720703125, 3339.01098632812, 
    3502.94213867188, 3635.50561523438, 3466.70971679688, 3395.76171875, 
    3546.62768554688, 3546.62768554688, 3575.19775390625, 3575.19775390625, 
    3572.06762695312, 3446.99755859375, 3348.94116210938, 3349.05639648438, 
    3349.05639648438, 3343.23461914062, 3228.00952148438, 3147.71850585938, 
    2904.17138671875, 2714.62939453125, 2736.48950195312, 2699.02294921875, 
    2881.1259765625, 3010.52856445312, 2970.4521484375, 3051.29931640625, 
    3051.29931640625, 3051.244140625, 3021.07861328125, 3045, 3045, 
    2983.88500976562, 2943.427734375, 2304.07641601562, 2616.2314453125, 
    2897.7509765625, 3047.69067382812, 3510, 3510, 3510, 2716.62109375, 
    2603.1279296875, 2816.537109375, 2949.45434570312, 2971.22338867188, 
    2939.18579101562, 2842.74340820312, 2810.67016601562, 3025, 3025, 
    2721.2265625, 2381.69677734375, 2470.71020507812, 2765.06225585938, 
    2855.17919921875, 2939.90014648438, 2884.30712890625, 2862.8037109375, 
    2963.712890625, 3130.3203125, 3516.470703125, 3692.12353515625, 
    3531.97314453125, 3387.2978515625, 3446.93090820312, 3424.07763671875, 
    3800.64697265625, 3721.27612304688, 3761.13208007812, 3920.50219726562, 
    3941.6953125, 3950.05541992188, 3950.05541992188, 3763.56225585938, 
    3939.931640625, 3558.76318359375, 3871.6240234375, 4162.765625, 
    4129.107421875, 4182.65625, 4227.9951171875, 4310.72021484375, 
    4356.388671875, 4457.82666015625, 4576.68310546875, 4690.13427734375, 
    4690.13427734375, 4667.8623046875, 4570.009765625, 4849.14208984375, 
    4827.2685546875, 4885.65576171875, 4852.14453125, 4975.10791015625, 
    4985.46142578125, 4944.6494140625, 4959.47216796875, 4904.38330078125, 
    4914.5048828125, 4971.3818359375, 4972.90283203125, 5008.20556640625, 
    4975.82275390625, 4977.5166015625, 4943.65234375, 4976.755859375, 
    4998.23095703125, 5035.5859375, 5046.68212890625, 5047.83837890625, 
    5077.17578125, 5039.34716796875, 4990.9970703125, 4999.01611328125, 
    4998.5732421875, 5020.4287109375, 5028.38037109375, 4964.11474609375, 
    4965.51123046875, 4937.31787109375, 4953.92626953125, 4904.818359375, 
    4941.56298828125, 4907.09814453125, 4875.078125, 4839.2421875, 
    4782.705078125, 4656.943359375, 4739.34423828125, 4319.45166015625, 
    4459.59375, 4615.48779296875, 4692.826171875, 4750.08984375, 
    4673.2255859375, 4660.21435546875, 4560.72314453125, 4568.916015625, 
    4481.76708984375, 4337.33056640625, 4289.94873046875, 4183.88037109375, 
    4137.67822265625, 4015.2578125, 3997.20092773438, 3950.80590820312, 
    3632.89575195312, 3804.048828125, 3744.37255859375, 3603.0517578125, 
    3323.19750976562, 2987.04248046875, 2801.13842773438, 1212.44763183594, 
    435.258392333984, 435.258392333984, 220, -0, -0, -0, -0, -0, -0, -0, 
    280.162628173828, 331.846557617188, 537.852905273438, 1866.45043945312, 
    2466.66776221529, 2917.91455078125, 3167.91186523438, 3576.54736328125, 
    3822.20263671875, 4036.1767578125, 4233.68017578125, 4301.0966796875, 
    4449.95947265625, 4579.47412109375, 4720.67724609375, 4586.53466796875, 
    4768.50390625, 4636.798828125, 4723.24755859375, 4745.84130859375, 
    4745.84130859375, 4632.63720703125, 4824.78759765625, 4815.43359375, 
    4872.39306640625, 4852.16650390625, 4845.57373046875, 4905.0400390625, 
    4942.34912109375, 4922.28076171875, 5022.64794921875, 4934.53759765625, 
    4963.48828125, 4965.28759765625, 5064.3525390625, 5119.44287109375, 
    5053.779296875, 4987.17041015625, 4986.81494140625, 5008.87548828125, 
    5044.97021484375, 5044.97021484375, 5008.80029296875, 5055.318359375, 
    5094.4638671875, 5078.6611328125, 5074.47509765625, 5126.494140625, 
    5133.36962890625, 5174.75537109375, 5168.23388671875, 5143.41858983545, 
    5199.63037109375, 5102.5517578125, 5160.0947265625, 5154.919921875, 
    5108.31689453125, 3971.59716796875, 2690.63012695312, 2180.771484375, 
    2319.5419921875, 2735.72607421875, 3548.60302734375, 3924.14428710938, 
    4743.66650390625, 4575.53466796875, 4868.7431640625, 4990.4599609375, 
    4837.79052734375, 4800.265625, 4786.35400390625, 4891.47509765625, 
    4808.75, 4806.26513671875, 5119.7158203125, 5024.9326171875, 
    5017.90380859375, 5061.62451171875, 4996.4150390625, 5017.462890625, 
    4955.86767578125, 5020.34130859375, 5035.150390625, 5100.94384765625, 
    5107.59228515625, 5089.7138671875, 5036.4521484375, 5023.9365234375, 
    4879.45849609375, 4651.51513671875, 4138.990234375, 4779.07571895829, 
    4779.07571895829, 4827.2451171875, 4907.0048828125, 4895.14404296875, 
    4828.54345703125, 4596.82763671875, 4374.1865234375, 4374.1865234375, 
    4345.4482421875, 4176.4365234375, 3798.85961914062, 3730.77465820312, 
    3125.84228515625, 3440.1884765625, 3440.1884765625, 3277.62377929688, 
    2932.72509765625, 3755.12182617188, 3721.27612304688, 3965.74243164062, 
    4017.48120117188, 3981.18310546875, 3968.43383789062, 3997.48803710938, 
    4108.87158203125, 4170.771484375, 3982.0068359375, 3644.18310546875, 
    3641.08642578125, 3770.43017578125, 3801.43530273438, 3638.69677734375, 
    3415.99951171875, 3218.10546875, 3140.28759765625, 3353.07592773438, 
    3398.39379882812, 3633.169921875, 3691.75805664062, 3461.22192382812, 
    3474.03149414062, 3471.80541992188, 3529.41967773438, 3534.16088867188, 
    3540.70361328125,
  3534.70043945312, 3481.70849609375, 3475, 3475, 3446.46752929688, 
    3502.26879882812, 3660.8447265625, 3675.1884765625, 3700.912109375, 
    3813.7666015625, 3774.5439453125, 3704.0361328125, 3603.716796875, 
    3303.56323242188, 2992.10473632812, 2933.13403320312, 2551.23657226562, 
    2326.11303710938, 2001.84252929688, 1567.82238769531, 1434.5869140625, 
    1467.74658203125, 2112.79638671875, 2949.28369140625, 3466.294921875, 
    3466.294921875, 3401.46875, 3134.26000976562, 3482.44384765625, 
    3897.27783203125, 3881.08447265625, 3531.7822265625, 3496.400390625, 
    3391.169921875, 3094.07934570312, 3072.72265625, 3046.62866210938, 
    3197.84790039062, 3481.31787109375, 3654.125, 3792.97119140625, 
    3923.21264648438, 3771.25805664062, 3881.84814453125, 3967.52685546875, 
    3895.60034179688, 3987.81420898438, 3987.81420898438, 3956.19970703125, 
    4136.6435546875, 4103.73095703125, 4065.89147763595, 4090.1767578125, 
    3945.43212890625, 4037.97827148438, 4037.97827148438, 3791.59765625, 
    3702.81420898438, 3665.96533203125, 3843.90307617188, 3755.5791015625, 
    3816.40551757812, 3840.17407226562, 3891.478515625, 3793.08959960938, 
    3823.30444335938, 3889.69018554688, 3888.28051757812, 3785.88623046875, 
    3661.90844726562, 3661.1064453125, 3490.23681640625, 3349.05639648438, 
    3349.05639648438, 3292.39697265625, 3178.56176757812, 3151.50244140625, 
    2495.36938476562, 2560.654296875, 2612.57495117188, 2668.67211914062, 
    2792.18530273438, 2843.8525390625, 2918.08227539062, 2900.88232421875, 
    2932.595703125, 2901.77807617188, 2723.22875976562, 2551.43994140625, 
    2410.37548828125, 1817.98132324219, 2065.32861328125, 2210.68432617188, 
    2901.19995117188, 2799.75561523438, 3045, 3517.0595703125, 
    3550.8974609375, 3326.45434570312, 3329.44946289062, 3403.98413085938, 
    3437.7177734375, 3458.841796875, 3264.52758789062, 3369.06176757812, 
    3167.97924804688, 3182.2880859375, 3012.39697265625, 3028.02465820312, 
    2945.68139648438, 2762.2265625, 2526.93237304688, 2415.71313476562, 
    2561.28100585938, 2611.58984375, 2721.0947265625, 2542.16870117188, 
    2758.41088867188, 2878.1884765625, 3155, 3155, 2956.3310546875, 
    2645.60961914062, 2732.62182617188, 2908.615234375, 3103.10913085938, 
    3109.59252929688, 3176.80932617188, 3402.10888671875, 3401.9287109375, 
    3670.79638671875, 3844.60668945312, 3764.67138671875, 3838.10717773438, 
    3848.990234375, 3850.25463867188, 4172.80908203125, 4216.53564453125, 
    4316.74658203125, 4290.94140625, 4531.1396484375, 4548.31982421875, 
    4528.240234375, 4660.01171875, 4690.13427734375, 4748.74072265625, 
    4665.6904296875, 4741.11767578125, 4741.11767578125, 4801.66162109375, 
    4886.46630859375, 4779.32958984375, 4983.1083984375, 5090.07080078125, 
    5125.7919921875, 5124.02587890625, 5055.99951171875, 5041.66748046875, 
    5040.34033203125, 5033.1552734375, 5040.650390625, 5006.814453125, 
    5043.0498046875, 5091.96484375, 5074.87744140625, 5133.27294921875, 
    5133.27294921875, 5117.6943359375, 5143.41858983545, 5190.8701171875, 
    5163.6865234375, 5171.80712890625, 5149.2109375, 5176.8642578125, 
    5090.40625, 5076.36767578125, 5079.162109375, 5056.99658203125, 
    5102.38818359375, 5066.734375, 5030.849609375, 5053.52685546875, 
    5085.44140625, 4932.20751953125, 4945.33740234375, 4937.9677734375, 
    4830.3408203125, 4691.521484375, 4720.32470703125, 4765.52587890625, 
    4761.83544921875, 4761.83544921875, 4620.365234375, 4764.5966796875, 
    4724.7158203125, 4695.2783203125, 4700.19775390625, 4610.6748046875, 
    4528.32666015625, 4438.287109375, 4437.05517578125, 4294.4716796875, 
    4204.57470703125, 4172.17138671875, 3983.87475585938, 3916.962890625, 
    3910.29467773438, 3848.8740234375, 3778.39111328125, 3797.74438476562, 
    3663.00341796875, 3453.52783203125, 3495.21630859375, 3349.67138671875, 
    2501.26806640625, 683.282409667969, 326.990295410156, 220, 220, 80, 80, 
    -0, -0, 190, 190, 180, 476.384185791016, 600.744689941406, 
    1724.38903808594, 2226.09448242188, 3550, 3550, 3550, 3532.23388671875, 
    3537.791015625, 3537.791015625, 3727.8359375, 4098.6865234375, 
    4307.44921875, 4516.45751953125, 4635.94287109375, 4688.30712890625, 
    4676.42578125, 4557.294921875, 4628.28955078125, 4575.333984375, 
    4768.2744140625, 4705.31689453125, 4749.2255859375, 4764.52197265625, 
    4750.103515625, 4900.3486328125, 4896.314453125, 4871.5888671875, 
    4847.93701171875, 4859.02392578125, 4922.97900390625, 4989.423828125, 
    4906.59716796875, 4944.16552734375, 4996.5859375, 5029.84130859375, 
    5076.1904296875, 5044.97021484375, 5044.97021484375, 5030.01416015625, 
    5055.318359375, 5068.337890625, 5068.337890625, 5172.52587890625, 
    5213.81591796875, 5198.6982421875, 5205.08984375, 5212.779296875, 
    5252.4072265625, 5311.78369140625, 5268.24853515625, 5164.6025390625, 
    5179.021484375, 5150.9931640625, 5223.8251953125, 5201.58056640625, 
    4482.05029296875, 4665.8837890625, 4643.927734375, 4894.326171875, 
    4914.28515625, 4988.45166015625, 4969.7099609375, 5076.15283203125, 
    5076.15283203125, 5013.81982421875, 5393.4189453125, 5426.2744140625, 
    5082.533203125, 5064.1201171875, 5095.03369140625, 5068.97119140625, 
    4891.05078125, 4982.1796875, 5050.69775390625, 5098.97509765625, 
    5046.2685546875, 5070.01904296875, 5052.57275390625, 5118.7724609375, 
    5121.87158203125, 5182.50732421875, 5143.671875, 5120.109375, 
    5127.8818359375, 5096.037109375, 5021.66455078125, 5029.62646484375, 
    5029.328125, 5006.61669921875, 5093.8173828125, 5003.611328125, 
    4978.0068359375, 4959.16943359375, 4853.76904296875, 4768.81494140625, 
    4834.9541015625, 4786.416015625, 4698.88330078125, 4485.712890625, 
    4195.7236328125, 4452.6240234375, 4697.87890625, 4734.15283203125, 
    4734.15283203125, 4734.15283203125, 4611.92724609375, 4724.9345703125, 
    4810.1923828125, 4880.88037109375, 4803.69921875, 4664.521484375, 
    4491.4521484375, 4300.05078125, 4377.75634765625, 4377.75634765625, 
    4114.47216796875, 4065.89147763595, 4146.974609375, 3994.97314453125, 
    3947.86108398438, 3946.09228515625, 3737.8505859375, 3819.28955078125, 
    3783.98974609375, 3779.00854492188, 3779.96875, 3792.2294921875, 
    3822.46435546875, 3727.48999023438, 3790.3642578125, 3866.01953125, 
    3696.33325195312, 3650,
  3050, 3050, 3050, 3050, 3175, 3373.61108398438, 3660.8447265625, 
    3675.1884765625, 3700.912109375, 4004.27416992188, 3886.99145507812, 
    3922.15405273438, 3860.66064453125, 3678.96044921875, 3592.3388671875, 
    3736.25732421875, 3816.79614257812, 3670.361328125, 3701.42114257812, 
    3701.42114257812, 3779.63623046875, 3812.810546875, 4166.6015625, 
    4223.896484375, 4237.86865234375, 4185.671875, 4246.87451171875, 
    4079.19458007812, 3908.83984375, 3850.837890625, 3985.67700195312, 
    4024.35717773438, 4024.35717773438, 4024.35717773438, 3999.61645507812, 
    3960.64501953125, 3945.35229492188, 4033.60546875, 4112.21923828125, 
    4105.087890625, 4098.291015625, 4149.984375, 4198.3896484375, 
    4204.9052734375, 4202.767578125, 4196.79931640625, 4196.88232421875, 
    4236.54296875, 4267.48681640625, 4310.23388671875, 4408.81298828125, 
    4408.81298828125, 4406.1533203125, 4509.51025390625, 4425.998046875, 
    4201.79931640625, 4080.48291015625, 3954.83715820312, 3748.3408203125, 
    3783.06860351562, 4098.87158203125, 4126.74560546875, 4122.98681640625, 
    4097.32861328125, 4048.68408203125, 4028.36547851562, 4028.36547851562, 
    4002.8232421875, 3896.81860351562, 3908.58911132812, 3445.78515625, 
    3575.81518554688, 3287.6259765625, 3038.78051757812, 2907.17407226562, 
    2907.17407226562, 2289.93530273438, 2137.46923828125, 2136.349609375, 
    2411.32763671875, 2639.22583007812, 2854.0498046875, 2804.9892578125, 
    2598.33178710938, 2617.50244140625, 2691.68139648438, 2582.12133789062, 
    2415.27001953125, 1899.31335449219, 3275, 3275, 3642.75756835938, 
    3937.3916015625, 4202.2783203125, 4157.69091796875, 3980.29174804688, 
    3780.27563476562, 3787.87133789062, 3686.4443359375, 3794.54125976562, 
    3963.91723632812, 3756.06176757812, 4054.703125, 3894.13818359375, 
    3786.607421875, 3641.09106445312, 3545.134765625, 3337.35717773438, 
    3325.44555664062, 3310.45336914062, 3020.16943359375, 2878.17626953125, 
    2758.41088867188, 2622.5537109375, 2576.84765625, 2707.83081054688, 
    2721.9150390625, 2483.78295898438, 2723.68920898438, 3155, 3155, 
    2924.68872070312, 2853.15625, 2610.53393554688, 2727.17407226562, 
    2835.11596679688, 2924.74462890625, 3109.10693359375, 3165.23022460938, 
    3262.60400390625, 3465.41748046875, 3510.70288085938, 3580.04760742188, 
    3670.37426757812, 3837.63940429688, 3858.27075195312, 4039.52465820312, 
    4031.60278320312, 4166.396484375, 4284.96142578125, 4487.001953125, 
    4529.42822265625, 4634.55029296875, 4660.01171875, 4676.13818359375, 
    4684.203125, 4765.93408203125, 4741.11767578125, 4741.11767578125, 
    4822.849609375, 4822.4873046875, 4879.28955078125, 4837.775390625, 
    5015.5625, 5115.58642578125, 5128.224609375, 5122.9130859375, 
    5052.32958984375, 5015.4267578125, 4996.36669921875, 4926.47509765625, 
    4971.36962890625, 5021.33349609375, 5089.53369140625, 5074.87744140625, 
    5133.27294921875, 5133.27294921875, 5151.88818359375, 5143.41858983545, 
    5176.1181640625, 5201.21728515625, 5181.13134765625, 5146.7685546875, 
    5154.05224609375, 5090.40625, 5076.36767578125, 5065.26416015625, 
    5013.23046875, 4893.46875, 4979.7724609375, 4911.59326171875, 
    5011.033203125, 5080.052734375, 5077.7001953125, 5036.07958984375, 
    4983.5849609375, 4888.34765625, 4825.5751953125, 4793.19580078125, 
    4750.4482421875, 4779.14501953125, 4799.640625, 4821.10400390625, 
    4849.9208984375, 4792.1572265625, 4780.49609375, 4763.16650390625, 
    4703.70263671875, 4650.65771484375, 4695.8984375, 4725.287109375, 
    4612.6943359375, 4563.14599609375, 4481.2158203125, 4386.60498046875, 
    4231.1865234375, 4267, 4184.23779296875, 4052.46899414062, 
    4052.46899414062, 4049.76245117188, 3883.12231445312, 3663.15258789062, 
    3540.97021484375, 3328.37548828125, 3350.51000976562, 3350.51000976562, 
    1228.63745117188, 880, 880, 880, 770, 770, 481.298400878906, 475, 475, 
    610.520874023438, 610.520874023438, 1724.38903808594, 3034.85888671875, 
    3034.85888671875, 3356.87109375, 3291.74389648438, 3203.79443359375, 
    2980.28662109375, 2301.75390625, 2034.35998535156, 2683.03491210938, 
    3419.59448242188, 3466.13061523438, 3258.92407226562, 3732.20385742188, 
    4705.9150390625, 4557.294921875, 4397.83349609375, 4091.8759765625, 
    4395.482421875, 4440.3671875, 4419.18185522252, 4331.40087890625, 
    4310.83740234375, 4763.2119140625, 4765.78564453125, 4765.78564453125, 
    4818.7646484375, 4851.21484375, 4590.25732421875, 4847.6796875, 
    4910.533203125, 4779.07571895829, 4749.24951171875, 5038.3759765625, 
    4952.35498046875, 4962.17236328125, 5030.01416015625, 5030.01416015625, 
    4891.1923828125, 5068.337890625, 5115.55615234375, 5222.63134765625, 
    5165.7822265625, 5277.24365234375, 5156.86328125, 5228.2939453125, 
    5220.94384765625, 5203.39892578125, 5276.4775390625, 5306.3486328125, 
    5354.73828125, 5330.67626953125, 5347.16943359375, 5376.43505859375, 
    5422.54833984375, 5342.08642578125, 5469.08740234375, 5271.5078125, 
    5228.34228515625, 5183.4736328125, 5094.71044921875, 5112.515625, 
    5090.17138671875, 5013.81982421875, 5428.28466796875, 5335.92578125, 
    5064.81689453125, 4983.35986328125, 5044.03564453125, 5076.0625, 
    5109.013671875, 5077.568359375, 5050, 5094.24560546875, 5112.19921875, 
    5131.6669921875, 5131.6669921875, 5129.74462890625, 5121.87158203125, 
    5143.41858983545, 5177.44677734375, 5168.04736328125, 5150.03271484375, 
    5116.1533203125, 5115.2568359375, 5119.845703125, 5107.2060546875, 
    5112.6318359375, 5095.4599609375, 5092.62841796875, 5076.00439453125, 
    5067.6591796875, 5044.8544921875, 5056.232421875, 5053.31396484375, 
    4978.15673828125, 4867.75830078125, 4731.998046875, 4709.958984375, 
    4786.34326171875, 4967.96630859375, 5031.876953125, 5008.53857421875, 
    5029.77978515625, 5041.12646484375, 5047.541015625, 5025.0830078125, 
    4928.8369140625, 4834.13916015625, 4739.4482421875, 4634.7783203125, 
    4539.8076171875, 4548.55712890625, 4557.24755859375, 4458.390625, 
    4332.64404296875, 4346.00439453125, 4335.45654296875, 4375.8984375, 
    4368.1845703125, 4270.2802734375, 4121.8212890625, 4045.22143554688, 
    4045.22143554688, 4016.95849609375, 4018.81372070312, 3909.19995117188, 
    3915.76635742188, 3940.30200195312, 3909.66333007812, 3696.33325195312, 
    3050,
  3050, 3050, 3050, 3050, 3050, 3170.06201171875, 3604.890625, 
    3764.8779296875, 4040.02758789062, 4082.14770507812, 4147.66455078125, 
    4199.8759765625, 4163.42041015625, 4173.02587890625, 4176.86572265625, 
    4124.24072265625, 4264.7509765625, 4390.8212890625, 4348.5810546875, 
    4391.33837890625, 4561.544921875, 4518.2392578125, 4519.69921875, 
    4510.0009765625, 4419.18185522252, 4185.671875, 4267.63037109375, 
    4267.63037109375, 4237.2626953125, 4185.712890625, 4176.98828125, 
    4161.32568359375, 4335.63671875, 4338.95751953125, 4297.7705078125, 
    4264.18408203125, 4304.5107421875, 4266.630859375, 4234.923828125, 
    4192.47509765625, 4217.74609375, 4304.01513671875, 4393.36572265625, 
    4404.236328125, 4365.98193359375, 4371.77783203125, 4419.18185522252, 
    4419.18185522252, 4458.275390625, 4499.232421875, 4556.03173828125, 
    4551.06494140625, 4514.3056640625, 4506.24951171875, 4518.7490234375, 
    4384.41064453125, 4301.35205078125, 4312.642578125, 4317.4619140625, 
    4289.14501953125, 4261.0205078125, 4308.568359375, 4247.98779296875, 
    4268.16064453125, 4209.947265625, 4028.36547851562, 4028.36547851562, 
    3983.77783203125, 3843.28442382812, 3887.46142578125, 3532.96313476562, 
    3243.1279296875, 2885.5810546875, 2746.57446289062, 2826.8115234375, 
    2780.72290039062, 2731.42211914062, 2602.86303710938, 2478.28759765625, 
    2323.58911132812, 2278.22216796875, 2651.26513671875, 2916.82788085938, 
    2893.29028320312, 2649.8916015625, 2831.88793945312, 2933.4619140625, 
    3400.6328125, 4154.7197265625, 4215.794921875, 3997.41040039062, 
    4522.154296875, 4517.234375, 4384.25341796875, 4391.68115234375, 
    4391.68115234375, 4348.9140625, 4387.86865234375, 4207.333984375, 
    4272.43408203125, 4172.9443359375, 4017.73120117188, 3934.533203125, 
    3922.73999023438, 3922.73999023438, 3886.70629882812, 3749.28076171875, 
    3851.51049804688, 3851.51049804688, 3548.45581054688, 3445.5419921875, 
    3218.02001953125, 3251.84692382812, 3465.91723632812, 3496.26342773438, 
    3660.91088867188, 3571.861328125, 3445.10815429688, 3493.0751953125, 
    3596.66015625, 3122.25927734375, 3275.89892578125, 3122.61254882812, 
    2834.48852539062, 2912.12768554688, 2811.63500976562, 2729.36962890625, 
    2766.59301757812, 2975.9990234375, 3125.26098632812, 3264.53686523438, 
    3468.13647460938, 3409.00732421875, 3538.9765625, 3669.55053710938, 
    3672.49267578125, 3904.8994140625, 3893.59204101562, 4002.87377929688, 
    4015.38330078125, 4015.38330078125, 4065.89147763595, 4307.08154296875, 
    4368.79443359375, 4387.84130859375, 4387.84130859375, 4660.10107421875, 
    4593.20751953125, 4699.40380859375, 4590.59814453125, 4522.61083984375, 
    4648.17578125, 4446.3466796875, 5015.5625, 5058.1533203125, 
    5073.669921875, 5074.2373046875, 5052.32958984375, 4993.4716796875, 
    4937.11328125, 4955.27490234375, 4967.048828125, 5079.833984375, 
    5042.2216796875, 5068.22705078125, 5044.53076171875, 5073.3544921875, 
    5181.7763671875, 5203.208984375, 5206.48291015625, 5193.966796875, 
    5082.23486328125, 5066.0888671875, 5051.88427734375, 5040.36328125, 
    4984.0888671875, 5086.8798828125, 5045.48876953125, 4952.94775390625, 
    5119.97998046875, 5119.97998046875, 5011.033203125, 5011.033203125, 
    5001.36572265625, 4992.017578125, 4908.27587890625, 4952.619140625, 
    4938.486328125, 4921.8271484375, 4842.482421875, 4876.04443359375, 
    4834.703125, 4826.5791015625, 4824.240234375, 4856.90576171875, 
    4790.099609375, 4732.5244140625, 4818.0322265625, 4847.556640625, 
    4878.1279296875, 4965.287109375, 4762.0498046875, 4762.0498046875, 
    4682.2314453125, 4537.8896484375, 4368.06884765625, 4324.2998046875, 
    4302.9580078125, 4296.64306640625, 4182.20703125, 4166.5732421875, 
    4029.64477539062, 3663.15258789062, 3540.97021484375, 3327.42211914062, 
    3544.53759765625, 3462.69067382812, 3476.50537109375, 4049.44018554688, 
    3721.27612304688, 2859.83447265625, 1850, 1056.06994628906, 985, 880, 
    880, 880, 880, 1529.11157226562, 3034.85888671875, 3034.85888671875, 
    3023.35913085938, 2550, 370.154968261719, 339.603088378906, 
    341.592956542969, 413.953002929688, 829.461669921875, 1101.54602050781, 
    3024.88842773438, 3024.88842773438, 2758.68920898438, 2791.4296875, 
    2791.4296875, 2168.89331054688, 2747.87475585938, 2747.87475585938, 
    3309.4775390625, 3219.97680664062, 3721.27612304688, 3825.82177734375, 
    4003.7197265625, 4003.7197265625, 4233.265625, 4279.06640625, 
    4242.08349609375, 4150, 4265.2431640625, 4265.2431640625, 4338.0234375, 
    4335.05126953125, 4534.20166015625, 4701.0634765625, 4514.89306640625, 
    4779.07571895829, 4826.197265625, 4779.07571895829, 4701.73779296875, 
    4708.5185546875, 4893.314453125, 5106.59521484375, 5124.92431640625, 
    4952.802734375, 5250.19287109375, 5236.07373046875, 5273.49609375, 
    5229.95458984375, 5294.44580078125, 5355.30126953125, 5392.564453125, 
    5395.818359375, 5403.0869140625, 5362.20166015625, 5352.087890625, 
    5336.31982421875, 5297.2421875, 5259.96337890625, 5272.81884765625, 
    5120.76171875, 5009.29931640625, 5015, 5015, 5015, 5280.00244140625, 
    5210.05615234375, 5186.44140625, 5050, 5010.939453125, 5043.53125, 
    5066.625, 5180.89697265625, 5301.82568359375, 5202.2431640625, 
    5152.98974609375, 5131.6669921875, 5173.2119140625, 5183.89111328125, 
    5218.333984375, 5234.6826171875, 5234.12841796875, 5217.8505859375, 
    5185.3505859375, 5190.7255859375, 5183.94482421875, 5173.0537109375, 
    5205.14892578125, 5233.52685546875, 5253.9990234375, 5229.84423828125, 
    5219.427734375, 5226.681640625, 5224.25732421875, 5211.0498046875, 
    5199.42626953125, 5162.49365234375, 5143.41858983545, 5143.41858983545, 
    5143.41858983545, 5171.306640625, 5194.833984375, 5200.8115234375, 
    5199.888671875, 5163.6943359375, 5117.2734375, 5065.1171875, 
    5030.1611328125, 4966.310546875, 4876.357421875, 4786.552734375, 
    4702.1357421875, 4703.642578125, 4441.78515625, 4458.51708984375, 
    4469.76904296875, 4406.64111328125, 4447.69482421875, 4422.78857421875, 
    4368.1845703125, 4387.888671875, 4201.47021484375, 4089.53979492188, 
    4192.4013671875, 4016.95849609375, 4039.1279296875, 4035.40185546875, 
    3862.15502929688, 3781.87548828125, 3536.60888671875, 3198.5361328125, 
    3050,
  2000, 1594.33801269531, 1628.88159179688, 1522.02001953125, 
    2467.3408203125, 3544.14697265625, 4011.6982421875, 4370.16259765625, 
    4370.16259765625, 4345.05615234375, 4326.81640625, 4303.32177734375, 
    4268.388671875, 4268.388671875, 4230.22705078125, 4388.15234375, 
    4419.18185522252, 4419.18185522252, 4424.0439453125, 4526.65380859375, 
    4647.91455078125, 4562.87744140625, 4467.00927734375, 4419.18185522252, 
    4455.34716796875, 4147.572265625, 4267.63037109375, 4269.5107421875, 
    4285.94189453125, 4397.40771484375, 4330.61328125, 4266.765625, 
    4320.13623046875, 4408.1484375, 4471.69287109375, 4518.60791015625, 
    4463.9736328125, 4375.26806640625, 4382.947265625, 4360.58251953125, 
    4408.44921875, 4376.1484375, 4393.521484375, 4505.22119140625, 
    4559.7822265625, 4511.64599609375, 4550, 4536.2041015625, 
    4552.4501953125, 4614.2021484375, 4624.09423828125, 4639.2392578125, 
    4606.234375, 4631.11083984375, 4623.47509765625, 4548.22314453125, 
    4459.47509765625, 4474.97705078125, 4407.61767578125, 4303.33740234375, 
    4276.4453125, 4221.1259765625, 4305.2470703125, 4274.72509765625, 
    4252.4609375, 4028.36547851562, 3803.7900390625, 3457.8134765625, 
    3481.04614257812, 3481.04614257812, 3143.0263671875, 3037.98583984375, 
    2930.48559570312, 2479.57250976562, 2860.69384765625, 2962.50122070312, 
    2962.50122070312, 2828.98706054688, 2765.22583007812, 2635.4482421875, 
    3118.52075195312, 3206.1884765625, 3507.48022460938, 3611.4619140625, 
    3468.05615234375, 3698.07641601562, 4223.1171875, 4419.18185522252, 
    4635.14794921875, 4643.41455078125, 4795.64599609375, 4779.07571895829, 
    4667.60693359375, 4681.35302734375, 4391.68115234375, 4391.68115234375, 
    4348.9140625, 4677.923828125, 4627.154296875, 4285.24951171875, 
    4232.4111328125, 4154.57275390625, 4141.01953125, 4132.96826171875, 
    4090.10815429688, 4077.73046875, 3930.24194335938, 4231.6005859375, 
    4102.6240234375, 3911.53759765625, 4072.498046875, 4327.60400390625, 
    4065.89147763595, 4115.689453125, 4244.4990234375, 3975.31079101562, 
    3733.85034179688, 3906.78295898438, 3948.55810546875, 3735.85571289062, 
    3539.0673828125, 3542.37817382812, 3431.25610351562, 3368.15625, 
    3276.59985351562, 3088.21484375, 2835.59423828125, 2575.7900390625, 
    2784.20776367188, 2892.13452148438, 3102.58178710938, 3220.32397460938, 
    3304.57861328125, 3345.8740234375, 3417.83666992188, 3465.5322265625, 
    3624.38696289062, 3609.38598632812, 3601.4853515625, 3696.123046875, 
    3949.6923828125, 4065.89147763595, 4257.61572265625, 4192.021484375, 
    4371.435546875, 4387.17333984375, 4369.59033203125, 4369.59033203125, 
    4302.4365234375, 4231.287109375, 4011.2822265625, 4285.4892578125, 
    4406.8740234375, 4900.42919921875, 5102.31201171875, 4697.5419921875, 
    4558.73095703125, 4730.7529296875, 4730.7529296875, 4721.7021484375, 
    4753.47705078125, 4896.64794921875, 4929.60498046875, 5044.0185546875, 
    5103.97412109375, 5044.53076171875, 5132.78369140625, 5132.78369140625, 
    5193.26611328125, 5174.3662109375, 5143.41858983545, 5082.23486328125, 
    4809.734375, 5040.36328125, 5040.36328125, 4974.76904296875, 
    5087.1494140625, 5045.48876953125, 4952.94775390625, 5124.18994140625, 
    5119.97998046875, 4817.68505859375, 4814.34326171875, 5025.2939453125, 
    5054.1611328125, 4972.91650390625, 4953.3349609375, 4871.798828125, 
    5057.0078125, 4895.431640625, 4895.431640625, 4902.544921875, 
    4933.98876953125, 4935.77978515625, 4859.703125, 4929.2392578125, 
    4909.56201171875, 4977.11572265625, 4944.46826171875, 4981.5146484375, 
    4974.3271484375, 4946.74658203125, 4862.24462890625, 4692.53466796875, 
    4571.15380859375, 4368.06884765625, 4324.2998046875, 4297.17919921875, 
    4221.89794921875, 4253.30224609375, 4185.12109375, 3895.2119140625, 
    3376.40014648438, 3525, 3525, 3525, 3646.32543945312, 3897.06958007812, 
    3721.27612304688, 3743.68359375, 3317.90063476562, 3552.767578125, 
    3578.56860351562, 3578.06225585938, 3525.779296875, 2550, 
    1924.61999511719, 1885, 2580.16748046875, 2580.16748046875, 
    2077.14794921875, 2077.14794921875, 1967.59631347656, 1750, 1750, 
    1831.79638671875, 3036.67138671875, 3036.67138671875, 2580.4814453125, 
    2388.53979492188, 2252.35815429688, 2252.35815429688, 1915.37292480469, 
    1634.728515625, 2057.29809570312, 2746.18823242188, 2746.18823242188, 
    2550, 2550, 2337.55517578125, 2257.193359375, 2434.13305664062, 
    1892.4345703125, 3960.05249023438, 4036.35888671875, 4150, 4150, 4150, 
    4150, 3278.36328125, 3278.36328125, 3130.02563476562, 3479.54174804688, 
    3935.43481445312, 4044.35083007812, 4150, 4561.33349609375, 
    4682.845703125, 4631.0478515625, 4621.13525390625, 4849.90283203125, 
    4949.99462890625, 4952.802734375, 5164.234375, 5236.265625, 
    5105.8095703125, 5235.8369140625, 5281.181640625, 5343.0703125, 
    5295.10400390625, 5340.88671875, 5333.958984375, 5328.4697265625, 
    5355.3427734375, 5327.287109375, 5316.5087890625, 5332.552734375, 
    5287.7900390625, 5133.12255859375, 5133.12255859375, 5130.9033203125, 
    5060.54541015625, 5058.890625, 5216.0458984375, 5342.728515625, 
    5187.5888671875, 5123.591796875, 5013.138671875, 5050, 5066.625, 
    5143.41858983545, 5245.74462890625, 5187.10205078125, 5350.61083984375, 
    5054.4248046875, 5264.89697265625, 5255.86572265625, 5261.6630859375, 
    5278.25830078125, 5277.9140625, 5257.23681640625, 5261.1494140625, 
    5235.3330078125, 5230.80615234375, 5272.48095703125, 5292.46533203125, 
    5281.42822265625, 5274.498046875, 5255.478515625, 5290.4892578125, 
    5288.29150390625, 5258.07763671875, 5250.873046875, 5252.13330078125, 
    5280.7431640625, 5275.79296875, 5275.021484375, 5274.93408203125, 
    5286.859375, 5273.4169921875, 5253.48779296875, 5242.248046875, 
    5212.14892578125, 5176.27490234375, 5131.76513671875, 5098.92724609375, 
    5025.64404296875, 4941.14306640625, 4921.1826171875, 4831.55712890625, 
    4732.2392578125, 4692.0703125, 4740.47412109375, 4608.5439453125, 
    4560.38134765625, 4580.68017578125, 4511.748046875, 4419.18185522252, 
    4373.31103515625, 4365.8017578125, 4332.09423828125, 4358.41748046875, 
    3751.67309570312, 3434.49169921875, 3137.70751953125, 2478.68994140625, 
    2972.384765625, 2972.384765625, 2876.18579101562, 2471.28540039062,
  1941.58776855469, 1594.33801269531, 1390.70678710938, 1552.92590332031, 
    2350.53149414062, 4231.9189453125, 4568.06689453125, 4689.625, 
    4604.7802734375, 4511.79638671875, 4590.6552734375, 4496.57958984375, 
    4498.79833984375, 4525.97265625, 4438.33935546875, 4388.15234375, 
    4452.08251953125, 4490.7744140625, 4509.091796875, 4493.822265625, 
    4399.2421875, 4338.06982421875, 4391.310546875, 4616.712890625, 
    4419.18185522252, 4266.9384765625, 4319.23974609375, 4385.619140625, 
    4385.619140625, 4396.40625, 4396.40625, 4521.5830078125, 4551.0576171875, 
    4587.23583984375, 4549.35546875, 4568.75830078125, 4594.8046875, 
    4597.45068359375, 4551.65771484375, 4578.74951171875, 4503.341796875, 
    4556.9462890625, 4514.18212890625, 4548.05322265625, 4624.84912109375, 
    4652.9189453125, 4670.61767578125, 4692.69091796875, 4636.86962890625, 
    4721.994140625, 4674.65869140625, 4682.5703125, 4675.59814453125, 
    4656.23046875, 4678.892578125, 4705.2607421875, 4587.82275390625, 
    4506.22265625, 4350.94091796875, 4190.67333984375, 4132.9697265625, 
    4300.4140625, 4202.78662109375, 4041.234375, 3844.9248046875, 
    3815.34545898438, 3645.82373046875, 3163.98046875, 3180.6201171875, 
    3127.55297851562, 3145, 3145, 3145, 2860.69384765625, 2860.69384765625, 
    3575, 3575, 3575, 3575, 3795.29296875, 3801.59594726562, 3615, 
    4097.37939453125, 4190.09033203125, 4403.31982421875, 4403.31982421875, 
    4683.93115234375, 4814.8564453125, 5033.04150390625, 4958.359375, 
    5013.2783203125, 5077.73486328125, 4824.5615234375, 4891.09130859375, 
    4965.71630859375, 5029.009765625, 4888.232421875, 4910.60009765625, 
    5050.1142578125, 4634.33740234375, 4630.90625, 4514.369140625, 
    4620.025390625, 4525.79296875, 4690.07373046875, 4697.72802734375, 
    4432.22509765625, 4310.291015625, 4367.73583984375, 4376.93896484375, 
    4376.93896484375, 4256.984375, 4291.740234375, 4308.12353515625, 
    4188.662109375, 4363.27978515625, 4354.71240234375, 4280.72998046875, 
    4260.03515625, 4021.31225585938, 3812.49584960938, 3612.2734375, 
    3646.33325195312, 3552.86450195312, 3394.1845703125, 3160.83178710938, 
    3017.86791992188, 2719.8798828125, 2533.08666992188, 2708.38647460938, 
    2705.0947265625, 2919.095703125, 3094.59716796875, 3160.50170898438, 
    3278.34643554688, 3200.0078125, 3359.966796875, 3375, 3516.12890625, 
    3586.75170898438, 3921.58325195312, 3987.1103515625, 3885.86401367188, 
    4103.435546875, 4162.93701171875, 4122.31640625, 4127.51171875, 
    4195.248046875, 4266.3681640625, 4100.498046875, 4011.2822265625, 
    4218.5146484375, 4218.5146484375, 4325.3310546875, 4419.9833984375, 
    4585.099609375, 4536.89111328125, 4567.94970703125, 4607.208984375, 
    4612.59033203125, 4636.76513671875, 4748.8076171875, 5039.6484375, 
    4910.6533203125, 5013.3623046875, 5013.1513671875, 5132.78369140625, 
    5132.78369140625, 5177.08642578125, 5202.46142578125, 5249.4970703125, 
    4759.36474609375, 4759.48828125, 4779.07571895829, 4872.4345703125, 
    5089.78759765625, 4997.9384765625, 4735.50634765625, 4790.8154296875, 
    4877.60400390625, 4940.5947265625, 4830.6708984375, 4845.65673828125, 
    4631.30126953125, 4568.65625, 4710.6396484375, 4919.064453125, 
    5035.10009765625, 4848.87744140625, 4910.828125, 4895.431640625, 
    5000.76025390625, 4988.9208984375, 4968.82421875, 4968.82421875, 
    5050.373046875, 5071.52392578125, 5097.75927734375, 5097.97607421875, 
    4819.87353515625, 5084.96923828125, 5005.880859375, 4847.37646484375, 
    4791.07666015625, 4768.52490234375, 4597.2109375, 4489.49169921875, 
    4403.75146484375, 4365.68798828125, 3949.8935546875, 3950, 3850, 3600, 
    3525, 3525, 3600, 3646.32543945312, 3933.720703125, 3867.21606445312, 
    3892.08862304688, 3525, 3552.767578125, 3581.20483398438, 
    3578.06225585938, 3801.80688476562, 3844.11206054688, 3636.87475585938, 
    3543.73974609375, 3019.63916015625, 3184.68676757812, 3550.62915039062, 
    3550.62915039062, 3550, 3375, 3375, 3375, 3375, 3375, 3040.02856445312, 
    3050, 3050, 3050, 3050, 2064.40161132812, 1482.39965820312, 2336.8203125, 
    2336.8203125, 2550, 2550, 3004.9580078125, 2963.49365234375, 
    2200.19287109375, 1307.66967773438, 2060.6962890625, 2949.19799804688, 
    4184.1923828125, 4184.1923828125, 4150, 4177.7294921875, 4173.9912109375, 
    3529.67578125, 3334.57397460938, 2867.49169921875, 3396.56909179688, 
    3890.11474609375, 4150, 4286.7900390625, 4243.16357421875, 
    4321.1279296875, 4548.62548828125, 4602.5791015625, 4827.2822265625, 
    4880.16650390625, 5119.7978515625, 5119.7978515625, 5105.8095703125, 
    5123.3076171875, 5121.93798828125, 5410.3203125, 5317.45849609375, 
    5107.07958984375, 5040.26025390625, 5207.6162109375, 5174.2509765625, 
    5148.08349609375, 5143.41858983545, 5251.15478515625, 5148.92236328125, 
    5133.12255859375, 5133.12255859375, 5181.58544921875, 5163.25146484375, 
    5246.38232421875, 5223.39501953125, 5314.974609375, 5202.52734375, 
    5123.7421875, 5057.11083984375, 5004.9609375, 5014.0126953125, 
    5100.3603515625, 5185.8876953125, 5321.6728515625, 5311.27197265625, 
    5453.68701171875, 5159.75732421875, 5314.03271484375, 5357.73095703125, 
    5316.39306640625, 5306.265625, 5270.7236328125, 5321.80517578125, 
    5296.54052734375, 5263.99951171875, 5251.10986328125, 5303.20556640625, 
    5292.962890625, 5313.31689453125, 5317.7314453125, 5317.1318359375, 
    5290.2392578125, 5286.33154296875, 5276.84521484375, 5302.56201171875, 
    5303.46435546875, 5312.37158203125, 5324.31494140625, 5334.037109375, 
    5333.533203125, 5322.51904296875, 5264.216796875, 5263.44287109375, 
    5220.3916015625, 5189.90576171875, 5185.48291015625, 5121.3564453125, 
    5072.796875, 5010.3603515625, 4932.6005859375, 4881.38623046875, 
    4856.38134765625, 4811.611328125, 4917.71728515625, 4685.33837890625, 
    4598.13671875, 4421.4697265625, 4748.6240234375, 4554.46337890625, 
    4459.04248046875, 4404.82177734375, 4232.5078125, 4232.5078125, 
    4178.26953125, 2274.87158203125, 1606.931640625, 1343.12084960938, 
    1235.07263183594, 1238.69079589844, 1622.40209960938, 1938.71472167969,
  1697.12502302956, 1700, 2079.65625, 2952.94165039062, 4215.6416015625, 
    4505.0673828125, 4690.22119140625, 4740.2412109375, 4740.2412109375, 
    4757.69091796875, 4637.6669921875, 4539.5322265625, 4557.80419921875, 
    4448.8564453125, 4419.18185522252, 4388.15234375, 4073.34350585938, 
    4243.36865234375, 4285.92919921875, 4260.3974609375, 4234.78564453125, 
    4333.3916015625, 4391.310546875, 4586.34375, 4419.18185522252, 
    4314.08203125, 4378.5869140625, 4385.619140625, 4385.619140625, 
    4396.40625, 4396.40625, 4514.08154296875, 4588.74169921875, 
    4559.10546875, 4498.71826171875, 4537.02880859375, 4714.20849609375, 
    4609.21435546875, 4697.35595703125, 4691.3076171875, 4584.1640625, 
    4620.1025390625, 4632.43359375, 4621.56103515625, 4587.06201171875, 
    4605.783203125, 4668.99169921875, 4636.98291015625, 4681.03564453125, 
    4681.03564453125, 4677.404296875, 4684.1787109375, 4688.765625, 
    4646.7529296875, 4620.81689453125, 4615.00537109375, 4612.50048828125, 
    4479.19482421875, 4253.216796875, 4155, 4155, 4167.7255859375, 
    4065.89147763595, 3867.90502929688, 3589.60815429688, 3441.05224609375, 
    3300.783203125, 3163.98046875, 3145, 3145, 3145, 3146.10278320312, 
    3294.26171875, 3157.23754882812, 3327.763671875, 3575, 3575, 3575, 3575, 
    3921.60424804688, 3795.29296875, 3615, 4202.6376953125, 4468.818359375, 
    4468.818359375, 4926.25537109375, 4964.31787109375, 5107.1064453125, 
    5231.9638671875, 5234.02978515625, 5177.71044921875, 5213.33642578125, 
    5256.55859375, 5189.2509765625, 5172.06640625, 4966.69873046875, 
    4978.58544921875, 4982.63720703125, 4922.17578125, 4985.5400390625, 
    4779.07571895829, 4830.60791015625, 4700.4365234375, 4526.55615234375, 
    4733.234375, 4755.658203125, 4755.658203125, 4615.43310546875, 
    4367.73583984375, 4376.93896484375, 4464.8759765625, 4560.79736328125, 
    4328.869140625, 4381.77685546875, 4567.12890625, 4428.11376953125, 
    4354.71240234375, 4333.16748046875, 4304.2431640625, 4021.31225585938, 
    3970.5478515625, 3919.05908203125, 3726.44262695312, 3684.349609375, 
    3605.0771484375, 3371.78955078125, 3123.39965820312, 2917.2744140625, 
    3051.10107421875, 2927.40161132812, 2758.41088867188, 2669.32983398438, 
    2886.16918945312, 2986.00122070312, 3121.53125, 3322.05932617188, 
    3326.46826171875, 3375, 3571.36694335938, 3661.96850585938, 
    3795.43725585938, 3721.27612304688, 3699.71142578125, 3513.00122070312, 
    3689.98413085938, 3979.63525390625, 3979.63525390625, 3463.13745117188, 
    3550.25463867188, 3687.326171875, 3836.23486328125, 3896.49731445312, 
    4165, 4165, 4325, 4334.93359375, 4452.0732421875, 4431.5185546875, 
    4695.64453125, 4531.97509765625, 4519.09326171875, 4595.86181640625, 
    4690.599609375, 4753.59619140625, 4907.37646484375, 4947.1318359375, 
    5101.77490234375, 5101.77490234375, 4752.376953125, 4752.376953125, 
    4708.55810546875, 4759.36474609375, 4759.36474609375, 4733.1015625, 4650, 
    4691.47802734375, 4564.701171875, 4541.9453125, 4595.41162109375, 
    4889.18017578125, 4885.70068359375, 4769.0595703125, 4769.0595703125, 
    4560, 4560, 4560, 4735.04833984375, 4908.1982421875, 4876.2822265625, 
    4966.80419921875, 4881.6640625, 4915.3154296875, 4899.70068359375, 
    4986.24462890625, 5073.53564453125, 5073.53564453125, 5043.92431640625, 
    4687.4111328125, 4747.35205078125, 4867.66259765625, 4860.72705078125, 
    4949.1806640625, 4855.38916015625, 4810.6982421875, 4768.52490234375, 
    4675.72900390625, 4533.31494140625, 4338.099609375, 3970.4130859375, 
    3950, 3950, 3850, 3600, 4050, 4050, 4050, 4050, 4050, 3700, 3525, 
    3683.8251953125, 3598.37280273438, 3578.06225585938, 4125, 4125, 
    4123.32861328125, 4086.46044921875, 3960.26733398438, 3674.314453125, 
    3550, 3550.62915039062, 3550.62915039062, 3550, 3375, 3375, 3375, 3375, 
    3375, 3200, 3200, 3200, 3200, 3200, 3200, 3200, 3200, 3200, 3200, 3200, 
    3291.97583007812, 3099.16943359375, 3285.84326171875, 3101.02856445312, 
    1775, 2047.99548339844, 4184.1923828125, 4553.1025390625, 
    4553.1025390625, 4306.126953125, 4128.02490234375, 4289.9755859375, 
    4294.0927734375, 3835.779296875, 3502.748046875, 3308.32397460938, 
    4203.171875, 4153.26708984375, 4150, 4252.5966796875, 4178.6435546875, 
    4268.50830078125, 4286.36376953125, 4535.1103515625, 4511.67138671875, 
    4509.2529296875, 4375.7314453125, 4698.31298828125, 4449.7626953125, 
    4550, 4550, 4614.61328125, 4515.48486328125, 4824.654296875, 
    5087.08203125, 5087.08203125, 5072.451171875, 5072.451171875, 
    4752.52001953125, 4606.6826171875, 4888.78515625, 5181.05078125, 
    5380.70751953125, 5500, 5500, 5411.02294921875, 5244.1171875, 
    5123.7421875, 4925.2919921875, 5028.29345703125, 4986.9443359375, 
    4906.173828125, 5008.75439453125, 5257.9697265625, 5365.28466796875, 
    5174.33544921875, 5292.4755859375, 5411.0029296875, 5372.1376953125, 
    5381.97216796875, 5406.4130859375, 5362.236328125, 5394.84033203125, 
    5348.4072265625, 5312.5927734375, 5343.9951171875, 5370.83056640625, 
    5344.20361328125, 5290.9208984375, 5263.29638671875, 5272.82958984375, 
    5124.89501953125, 5132.1923828125, 5286.23583984375, 5281.78857421875, 
    5333.009765625, 5340.955078125, 5323.65673828125, 5349.9990234375, 
    5365.97900390625, 5341.123046875, 5236.12060546875, 5244.0166015625, 
    5276.96630859375, 5225.92822265625, 5187.04052734375, 5104.83154296875, 
    5120.515625, 5066.12109375, 4963.95947265625, 4945.162109375, 
    4922.19873046875, 4914.11767578125, 4842.62841796875, 4682.01611328125, 
    4743.12353515625, 4206.31787109375, 4591.26318359375, 4433.96630859375, 
    4462.2763671875, 4404.82177734375, 4232.5078125, 4232.5078125, 
    4185.77490234375, 2970.927734375, 1995.65441894531, 1785, 1785, 1785, 
    1246.57482910156, 1370.53662109375,
  1877.96997070312, 2389.04760742188, 3734.07666015625, 4586.10302734375, 
    4677.95361328125, 4636.50439453125, 4719.64990234375, 4740.2412109375, 
    4740.2412109375, 4533.4072265625, 4503.83154296875, 4394.2353515625, 
    4169.0205078125, 4141.98974609375, 4134.0107421875, 4127.158203125, 
    4194.4677734375, 4276.01025390625, 4375.06787109375, 4269.80419921875, 
    4255.05126953125, 4264.84326171875, 4343.736328125, 4343.736328125, 
    4326.13427734375, 4314.08203125, 4371.83349609375, 4187.287109375, 
    4211.53759765625, 4300.90576171875, 4307.61865234375, 4466.0537109375, 
    4513.92626953125, 4496.8974609375, 4575.33349609375, 4629.40478515625, 
    4573.93115234375, 4678.5927734375, 4594.87646484375, 4594.87646484375, 
    4690.37353515625, 4726.7578125, 4796.203125, 4847.24853515625, 
    4755.64501953125, 4667.49658203125, 4666.91015625, 4690.16162109375, 
    4752.29345703125, 4742.38525390625, 4703.396484375, 4696.53369140625, 
    4579.291015625, 4505.3623046875, 4273.4755859375, 4247.5146484375, 
    4404.88134765625, 4404.1025390625, 4211.78125, 4002.96484375, 
    3957.28198242188, 3809.076171875, 3628.86840820312, 3521.57177734375, 
    3478.43505859375, 3148.56494140625, 3016.74389648438, 2900, 2900, 
    3222.45971679688, 3347.25146484375, 3239.41357421875, 3488.65356445312, 
    3508.33642578125, 3630.724609375, 3570, 3570, 3570, 2565, 
    3833.05639648438, 3738.34399414062, 3735.24560546875, 4202.6376953125, 
    4739.86083984375, 4642.091796875, 4988.580078125, 5094.15234375, 
    5023.79736328125, 5268.5390625, 5296.6328125, 5469.71728515625, 
    5336.68994140625, 5396.220703125, 5365.1357421875, 5427.20263671875, 
    5257.28173828125, 5112.93798828125, 5033.21875, 5085.08251953125, 
    5035.5048828125, 5063.74365234375, 4934.3310546875, 4893.75048828125, 
    4842.6708984375, 4733.234375, 4755.658203125, 4822.4892578125, 
    4782.11962890625, 4740.77001953125, 4678.3291015625, 4678.71728515625, 
    4464.8759765625, 4328.869140625, 4381.77685546875, 4454.00048828125, 
    4494.392578125, 4333.16748046875, 4344.99267578125, 4174.71142578125, 
    4113.732421875, 4197.0048828125, 4119.130859375, 3889.3623046875, 
    3743.205078125, 3695.48950195312, 3598.1455078125, 3311.78784179688, 
    3267.2080078125, 3172.43701171875, 3022.78930664062, 2877.220703125, 
    2612.88647460938, 2612.88647460938, 2597.33862304688, 2918.40112304688, 
    3086.51733398438, 3218.9306640625, 3375, 3610.2705078125, 
    3636.1533203125, 3703.07104492188, 3545.32666015625, 3088.70776367188, 
    3131.42895507812, 3282.26171875, 3491.24145507812, 3425.64916992188, 
    3457.25952148438, 3443.85083007812, 4165, 4165, 4160, 4165, 4165, 4265, 
    4265, 4350.94580078125, 4324.60107421875, 4357.51904296875, 
    4472.62939453125, 4595.1904296875, 4192.44873046875, 4740.923828125, 
    4690.599609375, 4583.9892578125, 4627.4482421875, 4717.99560546875, 
    4717.99560546875, 4454.92578125, 4386.31689453125, 4239.9560546875, 
    4500.78955078125, 4502.81689453125, 4597.3505859375, 4697.4951171875, 
    4583.27783203125, 4512.18408203125, 4419.18185522252, 4310, 
    4556.34814453125, 4572.8505859375, 4734.435546875, 4734.435546875, 
    4617.43359375, 4892.17919921875, 4930.18359375, 5143.431640625, 
    5208.873046875, 4711.51171875, 5102.96142578125, 5146.08740234375, 
    5143.41858983545, 5073.14599609375, 5199.60205078125, 5240.25244140625, 
    5087.2626953125, 4678.96240234375, 4940.82666015625, 4889.08740234375, 
    4735.3046875, 4735.3046875, 4655.27294921875, 4600.92529296875, 
    4603.4208984375, 4603.609375, 4472.69970703125, 4159.46728515625, 
    4090.07373046875, 3911.98852539062, 3975.03100585938, 3901.46313476562, 
    3850, 3699.66015625, 4050, 4050, 4050, 4050, 4050, 4050, 3700, 
    3768.1416015625, 4125, 4125, 4125, 4125, 4094.36352539062, 
    4366.60595703125, 4125, 4125, 3882.66748046875, 3939.751953125, 
    3667.19458007812, 3600, 3600, 3600, 3550, 3550, 3550, 3550, 
    3307.58520507812, 3200, 3200, 3303.42456054688, 3300, 3335.53344726562, 
    3365.79516601562, 3237.82299804688, 3301.57470703125, 3301.57470703125, 
    3223.44555664062, 3270.7392578125, 3346.783203125, 3070.06811523438, 
    1697.12502302956, 3505.80346679688, 4318.27587890625, 4553.1025390625, 
    4681.60009765625, 4506.19775390625, 4589.00634765625, 4690.27294921875, 
    4695.08203125, 4606.330078125, 4455.79443359375, 4250.21728515625, 
    4295.08642578125, 4295.08642578125, 4150, 4150, 3925.01684570312, 
    3784.47924804688, 3361.16918945312, 2859.39428710938, 3038.43969726562, 
    2864.85766601562, 3197.69384765625, 3324.37133789062, 3648.00854492188, 
    3769.13403320312, 3995.77587890625, 4042.03100585938, 4144.91796875, 
    4065.89147763595, 4148.11474609375, 4469.947265625, 4795.52001953125, 
    4878.80517578125, 4752.52001953125, 4933.77978515625, 5062.86669921875, 
    5160.34716796875, 5500, 5500, 5253.88525390625, 5467.69921875, 
    5414.05322265625, 5123.7421875, 5010.35888671875, 5048.27685546875, 4600, 
    4608.44140625, 4608.44140625, 4988.74951171875, 4988.74951171875, 
    5213.81787109375, 5299.001953125, 5327.94677734375, 5351.26025390625, 
    5395.638671875, 5427.203125, 5461.349609375, 5463.04736328125, 
    5466.0908203125, 5402.67578125, 5401.43212890625, 5393.97412109375, 
    5364.1826171875, 5143.41858983545, 5187.01318359375, 5277.1845703125, 
    5124.89501953125, 5132.1923828125, 5207.91259765625, 5190.10009765625, 
    5199.6845703125, 5154.35693359375, 5234.6328125, 5381.00439453125, 
    5382.30908203125, 5384.31103515625, 5330.22216796875, 5309.2119140625, 
    5350.9208984375, 5111.0068359375, 5111.0068359375, 5050.52734375, 
    4872.4287109375, 5008.8388671875, 4921.19287109375, 4869.93505859375, 
    4690.669921875, 4755.14208984375, 4708.30859375, 4617.1591796875, 
    4489.55322265625, 4206.31787109375, 4322.81103515625, 4322.81103515625, 
    3608.44140625, 2698.17407226562, 2650, 2693.47680664062, 
    2938.92358398438, 2938.92358398438, 2654.50317382812, 2486.55712890625, 
    2121.931640625, 2142.36596679688, 1699.68640136719, 1646.11193847656,
  3550, 4526.93017578125, 4482.50439453125, 4631.7802734375, 4545, 4545, 
    4545, 4531.82275390625, 4397.8330078125, 4117.041015625, 4040, 
    4044.13061523438, 4044.13061523438, 4127.18994140625, 4249.68408203125, 
    4355.455078125, 4243.9404296875, 4102.6494140625, 4044.91333007812, 
    4224.73291015625, 4151.5791015625, 4045, 4045, 4256.203125, 
    4242.5947265625, 4341.5966796875, 4199.94287109375, 4220.640625, 
    4130.7919921875, 4234.5439453125, 4369.6171875, 4471.49169921875, 
    4471.2568359375, 4435.1318359375, 4485.0810546875, 4495.92626953125, 
    4425.4384765625, 4444.0947265625, 4434.99462890625, 4553.291015625, 
    4625.2216796875, 4726.7578125, 4781.9521484375, 4784.822265625, 
    4755.64501953125, 4762.32568359375, 4666.91015625, 4676.22802734375, 
    4676.22802734375, 4640.728515625, 4581.48486328125, 4512.1416015625, 
    4419.19482421875, 4298.84765625, 4126.16357421875, 3876.0478515625, 
    3856.82299804688, 4045.40966796875, 4045.40966796875, 3915.59692382812, 
    3449.0791015625, 3526.7705078125, 3368.54736328125, 3188.68627929688, 
    3138.35498046875, 2793.33813476562, 2793.33813476562, 2902.12329101562, 
    3467.08276367188, 3434.54931640625, 3407.58422851562, 3501.21118164062, 
    3565.47143554688, 3576.0263671875, 3674.83911132812, 3689.65209960938, 
    3689.65209960938, 3689.65209960938, 1964.98132324219, 3974.48974609375, 
    3942.43017578125, 4065.89147763595, 4598.525390625, 4683.6962890625, 
    4683.6962890625, 4752.67822265625, 4751.73486328125, 5017.47265625, 
    5314.0654296875, 5178.51904296875, 5367.33203125, 5497.67529296875, 
    5441.68212890625, 5481.15576171875, 5346.58935546875, 5224.99560546875, 
    5005.990234375, 4994.98828125, 5028.16455078125, 5143.41858983545, 
    5143.41858983545, 5071.28857421875, 5001.8818359375, 4999.4619140625, 
    5028.7578125, 5018.1533203125, 5054.75927734375, 4970.634765625, 
    4863.18994140625, 4646.3369140625, 4610, 4610, 4610, 4516.80517578125, 
    4549.68115234375, 4442.77734375, 4333.86279296875, 4276.693359375, 
    4139.4296875, 4171.35546875, 4290.2060546875, 4218.8916015625, 
    4005.29321289062, 3754.93725585938, 3664.7197265625, 3568.3798828125, 
    3311.78784179688, 3351.68505859375, 3373.17724609375, 3364.58203125, 
    3186.43579101562, 2966.41723632812, 2846.07055664062, 2775.1005859375, 
    2716.30053710938, 2718.30395507812, 2909.83715820312, 3375, 3375, 
    2897.994140625, 2747.2890625, 2772.98120117188, 2896.99389648438, 
    3047.93041992188, 3237.74658203125, 3405.36450195312, 3445.42626953125, 
    3501.9345703125, 3628.6923828125, 4165, 4165, 4160, 4165, 4165, 
    4020.287109375, 3864.16381835938, 4245.1025390625, 4324.60107421875, 
    4324.60107421875, 4229.7294921875, 3872.4580078125, 3613.67407226562, 
    3585.92333984375, 3681.3603515625, 3793.18896484375, 3723.08178710938, 
    3825.16723632812, 4020.73071289062, 4043.43115234375, 4032.55834960938, 
    4065.89147763595, 4132.12255859375, 4133.96337890625, 4356.09228515625, 
    4354.3017578125, 4446.91650390625, 4494.0166015625, 4346.52734375, 
    4310.4208984375, 4367.42724609375, 4433.26416015625, 4655.14794921875, 
    4679.1025390625, 4617.43359375, 5033.3916015625, 5500, 5318.05908203125, 
    5155.64697265625, 5019.8056640625, 5102.96142578125, 5349.9814453125, 
    5343.46240234375, 5073.14599609375, 5359.31494140625, 5314.599609375, 
    4793.66943359375, 4926.58837890625, 4807.4560546875, 4817.2939453125, 
    4590.22314453125, 4662.8779296875, 4534.701171875, 4452.7685546875, 
    4319.154296875, 4278.091796875, 4271.53271484375, 4290.3466796875, 
    4075.83325195312, 3911.98852539062, 3548.2529296875, 3200, 3200, 3200, 
    3200, 3441.88842773438, 3441.88842773438, 4050.78149414062, 4125, 4125, 
    4125, 4125, 4125, 4125, 4125, 4125, 4125, 4125, 4125, 4120.375, 4120.375, 
    4025, 4025, 3692.87084960938, 4005.63891601562, 3798.15844726562, 3550, 
    3550, 3550, 3550, 3307.58520507812, 3200, 3200, 3356.53930664062, 3300, 
    3335.53344726562, 3367.7646484375, 3237.82299804688, 3327.00244140625, 
    3301.57470703125, 3300, 3310.10791015625, 2927.54760742188, 1850, 
    2932.38525390625, 4342.76171875, 4342.76171875, 4318.27587890625, 
    4419.18185522252, 4506.19775390625, 4683.330078125, 4690.27294921875, 
    4690.27294921875, 4677.587890625, 4462.5703125, 4404.1396484375, 
    4295.08642578125, 4295.08642578125, 4349.24560546875, 4201.61328125, 
    3987.07934570312, 3963.07666015625, 3687.86889648438, 3420.18872070312, 
    3065.78548661781, 2990.29028320312, 3044.33447265625, 3253.96899414062, 
    3547.00634765625, 3498.783203125, 3780.59985351562, 3914.7744140625, 
    4247.02197265625, 4169.416015625, 3901.078125, 4346.86328125, 
    4366.35595703125, 4349.79833984375, 4688.3427734375, 4933.77978515625, 
    5062.86669921875, 5192.00390625, 5344.171875, 5391.435546875, 
    5197.20849609375, 5176.6787109375, 5224.72802734375, 5122.666015625, 
    5017.89794921875, 4458.41064453125, 4408.76953125, 4300, 4300, 4300, 
    4300, 4952.12890625, 5219.90966796875, 5326.0400390625, 5408.47216796875, 
    5428.0810546875, 5453.32861328125, 5428.82080078125, 5464.54833984375, 
    5407.390625, 5331.6259765625, 5322.98681640625, 5354.63916015625, 
    5283.98876953125, 5086.84814453125, 4892.90185546875, 5117.47705078125, 
    5117.47705078125, 4929.0087890625, 4800.74560546875, 4925.046875, 
    4830.21630859375, 5003.99951171875, 5057.9814453125, 5143.41858983545, 
    5274.17578125, 5422.86767578125, 5421.7431640625, 5373.40283203125, 
    5169.8681640625, 5067.21630859375, 5059.22705078125, 4672.6318359375, 
    4595.9228515625, 4516.76904296875, 4848.9345703125, 4877.54736328125, 
    4690.669921875, 4708.30859375, 4708.30859375, 4617.1591796875, 
    4330.09033203125, 3393.71362304688, 2039.96069335938, 1288.07080078125, 
    1995.07397460938, 2942.54272460938, 2977.71118164062, 2650, 2650, 
    2654.50317382812, 2654.50317382812, 2581.70629882812, 2121.931640625, 
    2121.931640625, 1961.6015625, 2272.79223632812,
  3550, 4515.56884765625, 4637.8564453125, 4422.130859375, 4646.681640625, 
    4553.111328125, 4545.75830078125, 4419.18185522252, 4419.18185522252, 
    4433.79833984375, 4238.03857421875, 4128.82275390625, 4190.11669921875, 
    4225.95556640625, 4302.79833984375, 4300.2353515625, 3987.8828125, 
    3972.3232421875, 3934.42553710938, 3887.54858398438, 3939.84033203125, 
    3939.84033203125, 3885.767578125, 4098.46826171875, 4230.91064453125, 
    3950.46997070312, 3914.36401367188, 3974.31030273438, 3899.00512695312, 
    3863.67407226562, 4000.06176757812, 4212.39990234375, 4317.46240234375, 
    4517.79931640625, 4426.779296875, 4400.56005859375, 4400.56005859375, 
    4355.89306640625, 4354.16943359375, 4382.5673828125, 4505.40869140625, 
    4514.28466796875, 4590.02685546875, 4577.2861328125, 4600.63330078125, 
    4617.30322265625, 4620.64697265625, 4657.96923828125, 4431.79345703125, 
    4449.07421875, 4355.22119140625, 4248.5205078125, 4186.0732421875, 
    4050.76977539062, 3869.61303710938, 3820.947265625, 3964.15673828125, 
    3943.11401367188, 3929.40795898438, 3828.47924804688, 3617.4931640625, 
    3220.701171875, 3161.34887695312, 3080.72290039062, 2712.38671875, 
    2680.52416992188, 2539.16040039062, 3352.2275390625, 4055.78979492188, 
    3885.70434570312, 3703.72534179688, 3804.58154296875, 3838.2255859375, 
    3821.34448242188, 3924.98706054688, 4013.89184570312, 4049.48364257812, 
    4215, 4215, 4408.19091796875, 4381.42529296875, 4579.91357421875, 
    4598.525390625, 4683.6962890625, 4683.6962890625, 2289.51928710938, 
    1901.56579589844, 2365.0283203125, 3135.93505859375, 4645.5244140625, 
    5108.07958984375, 5447.4853515625, 5433.314453125, 5405.50146484375, 
    5291.9833984375, 5098.44921875, 5096.76416015625, 5117.05615234375, 
    5216.220703125, 5269.2294921875, 5220.08544921875, 5212.98046875, 
    5143.41858983545, 5223.3037109375, 5230.716796875, 5217.70751953125, 
    5004.14892578125, 4945.4580078125, 4865.482421875, 4633.34619140625, 
    4616.1826171875, 4682.4736328125, 4682.4736328125, 4607.7060546875, 
    4656.5888671875, 4656.5888671875, 4610, 4589.98974609375, 
    4277.79541015625, 4369.82861328125, 4167.10595703125, 4166.01416015625, 
    3977.13232421875, 3947.90258789062, 4039.20727539062, 3624.47534179688, 
    3402.05419921875, 3351.68505859375, 3482.70361328125, 3509.44677734375, 
    3405.45556640625, 3248.30444335938, 3155.61840820312, 3159.48559570312, 
    3193.5419921875, 3353.61987304688, 3353.61987304688, 3375, 3375, 
    2947.06884765625, 2747.2890625, 2594.94897460938, 2742.3896484375, 
    2904.81103515625, 3014.7529296875, 3091.66284179688, 3242.22680664062, 
    3279.6806640625, 3528.373046875, 4165, 4165, 3640.66430664062, 
    3534.35961914062, 3580, 3580, 3554.04907226562, 3387.2978515625, 
    2814.20043945312, 2481.9501953125, 2731.81396484375, 2963.93359375, 
    3071.15625, 3212.2099609375, 3509.19458007812, 3682.73754882812, 
    3726.78930664062, 3721.27612304688, 3621.35498046875, 3826.0078125, 
    3891.92626953125, 3966.095703125, 4031.11059570312, 3977.11376953125, 
    4065.89147763595, 4258.12060546875, 4370.3759765625, 4370.3759765625, 
    4346.52734375, 4406.04248046875, 4406.04248046875, 4350, 
    4576.37744140625, 4593.82177734375, 4556.5068359375, 5121.17236328125, 
    5451.572265625, 5367.4482421875, 5357.22900390625, 5019.8056640625, 
    5044.294921875, 5076.21875, 5076.21875, 4966.25634765625, 5105.068359375, 
    4838.73876953125, 4829.583984375, 5038.35302734375, 4927.0703125, 
    4701.71142578125, 4688.76416015625, 4472.5615234375, 4405.3466796875, 
    4152.958984375, 4088.04565429688, 3916.92749023438, 4151.18994140625, 
    4137.49462890625, 2413.990234375, 1652.36779785156, 985, 985, 985, 985, 
    985, 2366.50366210938, 3311.81713867188, 3834.92065429688, 4125, 4125, 
    4125, 4125, 4125, 4125, 3600, 3600, 2551.95458984375, 3723.84765625, 
    4125, 4233.43603515625, 4120.375, 4027.19506835938, 4025, 4025, 4025, 
    4025, 4025, 3525, 3525, 3525, 3199.13354492188, 3200, 3200, 
    2879.08129882812, 2725.419921875, 2725, 2725, 3225, 3225, 3550, 3550, 
    3550, 4125, 4849.5068359375, 4849.5068359375, 4694.77685546875, 
    4342.76171875, 4125, 4125.73681640625, 4263.09033203125, 
    4425.74365234375, 4425.74365234375, 4453.85986328125, 4467.9755859375, 
    4424.4169921875, 4079.07421875, 4043.802734375, 4055.58154296875, 
    4201.61328125, 4254.04736328125, 3987.07934570312, 3836.34375, 
    3687.86889648438, 3563.13061523438, 3368.19775390625, 2990.29028320312, 
    2888.10864257812, 3065.78548661781, 3188.9140625, 3214.62475585938, 
    3214.62475585938, 3547.29809570312, 3387.2978515625, 3414.869140625, 
    3120.6298828125, 3155.16528320312, 2985.43237304688, 3156.68725585938, 
    3665.69750976562, 4301.68505859375, 4328.8173828125, 4228.84033203125, 
    4950.974609375, 5109.19482421875, 5045.8271484375, 5102.82373046875, 
    5091.697265625, 4964.63525390625, 4634.7275390625, 4691.85986328125, 
    4210.96435546875, 3945.25122070312, 3891.1689453125, 3850, 3850, 
    4647.5546875, 4648.35009765625, 4648.35009765625, 5416.3037109375, 5500, 
    5484.330078125, 5473.68603515625, 5444.537109375, 5464.98779296875, 
    5381.78369140625, 5236.2177734375, 5201.271484375, 5179.92236328125, 
    4419.18185522252, 4009.42260742188, 4005, 4141.39501953125, 
    4352.615234375, 4222.28076171875, 4463.5205078125, 4554.87548828125, 
    4567.10009765625, 4621.2587890625, 4841.73046875, 5190.1650390625, 
    5285.517578125, 5206.88916015625, 5178.48388671875, 5223.6884765625, 
    5067.21630859375, 4985.87646484375, 4338.828125, 4338.828125, 
    4294.89697265625, 4650, 4663.22509765625, 4734.79541015625, 
    4612.4541015625, 4637.53271484375, 4501.212890625, 3835.56616210938, 
    2723.47973632812, 3194.9677734375, 4173.11669921875, 4270.99560546875, 
    4241.4619140625, 3439.33251953125, 3232.77294921875, 2975.90283203125, 
    2654.50317382812, 2654.50317382812, 2581.70629882812, 2120, 2120, 
    2373.54858398438, 2660.005859375,
  3590.15405273438, 3960.41040039062, 3805.20703125, 4293.30712890625, 
    4293.30712890625, 4585.46240234375, 4527.08349609375, 4545.92431640625, 
    4460.45263671875, 4470.35107421875, 4314.16455078125, 4202.7802734375, 
    4273.7509765625, 4263.51025390625, 4161.4560546875, 4014.80737304688, 
    3781.9296875, 3643.73876953125, 3763.51928710938, 3799.63696289062, 
    3653.96166992188, 3777.10205078125, 3979.8505859375, 3902.64599609375, 
    4042.13305664062, 3951.4521484375, 3970.39453125, 3826.01904296875, 
    3830.00756835938, 3833.08203125, 3733.60864257812, 3889.16552734375, 
    4042.65991210938, 4127.1337890625, 4175.41748046875, 4290.509765625, 
    4277.916015625, 4170.87451171875, 4230.8310546875, 4166.69287109375, 
    4295.52197265625, 4316.35595703125, 4368.79443359375, 4368.79443359375, 
    4612.12353515625, 4603.30859375, 4510.443359375, 4429.8876953125, 
    4358.64599609375, 4377.46728515625, 4222.89501953125, 4112.8466796875, 
    4065.89147763595, 3903.26586914062, 3849.43774414062, 3965.05004882812, 
    3836.943359375, 3739.046875, 3661.34521484375, 3661.34521484375, 
    3446.29125976562, 2871.68383789062, 2956.73828125, 2766.283203125, 
    2567.2421875, 2500.33276367188, 2969.37109375, 3600.00122070312, 
    3817.5703125, 3939.84033203125, 3654.03125, 3955.6455078125, 
    4019.34765625, 4133.0419921875, 4207.00244140625, 4089.07153320312, 
    4116.01025390625, 4215, 4215, 4381.42529296875, 4381.42529296875, 
    4578.56591796875, 4452.11474609375, 4574.8212890625, 1792.67895507812, 
    1393.26257324219, 1393.26257324219, 920.56396484375, 1043.94641113281, 
    1191.69055175781, 1750.31909179688, 3956.99096679688, 5001.76318359375, 
    5052.74853515625, 5052.74853515625, 4996.74560546875, 4834.0625, 
    4983.26171875, 5248.8515625, 5316.89453125, 5291.7841796875, 
    5373.26318359375, 5341.1328125, 5318.173828125, 5385.03125, 
    5278.13330078125, 5248.23681640625, 5216.4345703125, 5179.14013671875, 
    5063.4921875, 4883.77099609375, 4981.99658203125, 4936.37646484375, 
    4962.6513671875, 4885.1806640625, 4906.47265625, 4924.2255859375, 
    4578.591796875, 4487.9404296875, 4382.88720703125, 4340.537109375, 
    4152.16455078125, 4033.5361328125, 4033.5361328125, 3869.64770507812, 
    3611.85278320312, 3491.99682617188, 3656.17309570312, 3704.58959960938, 
    3704.58959960938, 3813.72509765625, 3928.95166015625, 3871.8427734375, 
    3536.18237304688, 3706.34008789062, 3611.21752929688, 3353.61987304688, 
    3375, 3375, 2947.06884765625, 2651.33618164062, 2411.27954101562, 
    2372.1611328125, 2589.32421875, 2636.68798828125, 2812.89135742188, 
    3130.80541992188, 3420.07055664062, 3496.01147460938, 4165, 4165, 
    3779.19311523438, 3535, 3580, 3580, 3183.22875976562, 3205.94604492188, 
    2950.69409179688, 2758.41088867188, 2701.65014648438, 2710.67993164062, 
    2710.67993164062, 2894.81494140625, 3093.06958007812, 3309.16259765625, 
    3334.61938476562, 3524.32177734375, 3520.47412109375, 3671.09545898438, 
    3827.5048828125, 3822.48950195312, 3920.53564453125, 3889.63647460938, 
    4112.271484375, 4094.94140625, 4065.89147763595, 4166.85302734375, 
    4284.89501953125, 4406.04248046875, 4408.77734375, 4382.587890625, 
    4486.1455078125, 4498.7021484375, 4504.052734375, 4851.87353515625, 
    5040.5390625, 5097.00537109375, 4934.560546875, 4503.5771484375, 
    4588.10302734375, 4515.96044921875, 4812.35693359375, 4977.54248046875, 
    5006.28369140625, 5001.4990234375, 4886.85107421875, 4845.2998046875, 
    4673.787109375, 4565.125, 4469.044921875, 4310.068359375, 
    4074.9892578125, 4065.89147763595, 3971.32373046875, 3916.92749023438, 
    2796.25146484375, 425.785466617812, 0, -0, -0, -0, -0, -0, -0, 40, 120, 
    190, 281.717864990234, 281.717864990234, 110, 140, 140, 140, 220, 
    1148.83056640625, 2551.95458984375, 3892.98779296875, 3904.90161132812, 
    3904.90161132812, 4025, 4025, 4025, 4025, 4025, 4052.013671875, 
    4014.40576171875, 3525, 3525, 3525, 2556.65234375, 2265.7470703125, 1350, 
    650, 485, 985, 2218.7001953125, 3225, 3225, 3550, 3550, 3550, 4125, 
    4849.5068359375, 4849.5068359375, 4694.77685546875, 4395.3642578125, 
    4294.005859375, 4209.09033203125, 4130.41455078125, 4008.73364257812, 
    4663.5537109375, 4556.5400390625, 4357.84033203125, 4126.7587890625, 
    4069.76879882812, 3992.22680664062, 3936.787109375, 3770.3798828125, 
    3858.82543945312, 3568.85620117188, 3237.26538085938, 3151.02612304688, 
    3243.62866210938, 2938.4169921875, 2568.20849609375, 2553.69311523438, 
    2588.76733398438, 2434.712890625, 2034.86694335938, 1999.78735351562, 
    2201.21484375, 2226.013671875, 2226.013671875, 1766, 2409.50659179688, 
    2786.55004882812, 2786.55004882812, 3360.95458984375, 3360.95458984375, 
    3469.73608398438, 4017.88012695312, 4140.1923828125, 4344.88671875, 
    4500.59375, 4728.61181640625, 4703.046875, 4419.18185522252, 
    4229.5537109375, 3930.09106445312, 3930.96044921875, 3655.61987304688, 
    3627.20727539062, 3627.20727539062, 3621.06811523438, 3792.17309570312, 
    3792.17309570312, 4711.14453125, 5014.60498046875, 5153.5771484375, 
    5364.90771484375, 5483.6787109375, 5399.5498046875, 5414.3505859375, 
    5424.77294921875, 5209.57373046875, 4917.49072265625, 4849.27294921875, 
    4320.3544921875, 3474.19140625, 3470, 3470, 3470, 3573.9423828125, 
    3816.19653320312, 4026.97338867188, 3957.1337890625, 4188.3505859375, 
    4441.962890625, 4441.962890625, 4185, 3255, 4185, 4185, 4335.55078125, 
    4528.40283203125, 4528.40283203125, 4365.5029296875, 4403.43359375, 4650, 
    4650, 4757, 4742.466796875, 4729.53076171875, 4705.02490234375, 
    4272.0361328125, 4419.18185522252, 4455.3173828125, 4400.93017578125, 
    4236.8212890625, 4065.89147763595, 3439.33251953125, 3232.77294921875, 
    2975.90283203125, 2004.93139648438, 1423.19921875, 1350.482421875, 2120, 
    2120, 2373.54858398438, 3399.16162109375,
  3445, 3445, 3494.9853515625, 4197.3994140625, 4375.63330078125, 
    4588.21337890625, 4578.66943359375, 4555.298828125, 4515.447265625, 
    4419.18185522252, 4314.16455078125, 4267.6806640625, 4180.4482421875, 
    4157.2041015625, 3965.33618164062, 3950.50073242188, 3991.37084960938, 
    3940.72680664062, 3822.19018554688, 3822.45556640625, 3674.68994140625, 
    3859.44653320312, 3854.29541015625, 3860.1279296875, 3765.24658203125, 
    3766.91772460938, 3827.99755859375, 3788.40307617188, 3859.10791015625, 
    3662.02661132812, 3633.376953125, 3758.98876953125, 3901.66821289062, 
    3845.91235351562, 4014.92138671875, 3953.92895507812, 4039.9345703125, 
    4027.48754882812, 4213.52392578125, 4109.2236328125, 4295.54345703125, 
    4380.5, 4368.79443359375, 4368.79443359375, 4479.7119140625, 
    4519.51611328125, 4519.4599609375, 4181.18798828125, 4207.84814453125, 
    4165.5830078125, 3898.2158203125, 3852.06640625, 3863.1865234375, 
    3959.29174804688, 3834.6494140625, 3695.08325195312, 3575.37841796875, 
    3556.1806640625, 3337.9501953125, 3337.9501953125, 3269.60131835938, 
    2937.1015625, 2935.6787109375, 2918.35571289062, 2909.9609375, 
    3023.6669921875, 4050, 4050, 4050, 4050, 4050, 4050, 4208.6943359375, 
    4182.05908203125, 4090.51123046875, 4225.95556640625, 4114.857421875, 
    4223.41552734375, 4295.2578125, 3612.51220703125, 3612.51220703125, 3615, 
    4241.5439453125, 4229.751953125, 3562.59448242188, 1335.96594238281, 
    1222.39440917969, 944.656433105469, 803.740539550781, 612.486755371094, 
    581.002014160156, 462.868927001953, 535.145141601562, 2226.69848632812, 
    4289.22607421875, 4970.45263671875, 4839.9423828125, 4839.44384765625, 
    4997.177734375, 5118.56884765625, 5315.3583984375, 5266.88427734375, 
    5403.7041015625, 5500, 5487.0234375, 5473.06982421875, 5499.9736328125, 
    5500, 5500, 5420.0888671875, 5193.42333984375, 5218.1376953125, 
    4981.3525390625, 4970.2060546875, 5008.9560546875, 4943.37939453125, 
    4906.47265625, 4666.98291015625, 4515, 4515, 4255.60595703125, 
    4229.83349609375, 4266.9296875, 4033.5361328125, 4036.5234375, 
    4036.5234375, 3982.15649414062, 4138.623046875, 4138.623046875, 
    4143.7255859375, 4166.3017578125, 4023.40844726562, 3983.45092773438, 
    3786.5458984375, 3797.30151367188, 3758.2197265625, 3465.5556640625, 
    3375, 3184.9755859375, 1999.78979492188, 2518.9091796875, 
    2908.98706054688, 3028.97338867188, 3034.56201171875, 3618.23364257812, 
    4202.3671875, 4202.3671875, 4187.4189453125, 4042.04907226562, 4165, 
    4165, 3858.42456054688, 3691.30078125, 3641.52758789062, 3610.6376953125, 
    3589.3837890625, 3356.58129882812, 3190.0986328125, 2971.33984375, 
    3037.24975585938, 2710.67993164062, 2710.67993164062, 2814.10083007812, 
    3187.35571289062, 3320.66015625, 3491.42431640625, 3503.7080078125, 
    3560.46850585938, 3616.31030273438, 3536.90942382812, 3747.83911132812, 
    3928.07495117188, 3927.94091796875, 4009.20947265625, 4077.16479492188, 
    4129.916015625, 4220.9921875, 4299.13623046875, 4256.60400390625, 
    4379.22265625, 4382.587890625, 4473.44970703125, 4461.5068359375, 
    4403.78076171875, 4667.52880859375, 4715.32470703125, 4802.2109375, 
    4922.35791015625, 4872.716796875, 4807.6328125, 4843.5517578125, 
    4990.05859375, 5007.78125, 5016.1494140625, 5035.99169921875, 
    4929.7958984375, 4675.939453125, 4689.390625, 4440.97607421875, 
    4345.24951171875, 4274.8525390625, 4094.412109375, 4007.66088867188, 
    4033.26904296875, 2176.08862304688, 819.895812988281, -0, -0, -0, -0, -0, 
    -0, 70, 90, 120, 150, 257.514770507812, 311.124694824219, 
    311.124694824219, 170, 140, 140, 426.629821777344, 1297.03967285156, 
    1592.55358886719, 2250.583984375, 2250.583984375, 1367.74340820312, 
    1296.98779296875, 1968.64721679688, 2324.66235351562, 3252.77490234375, 
    3252.77490234375, 2626.4794921875, 2626.4794921875, 1980.29516601562, 
    1915.23181152344, 1450, 1450, 2177.31420898438, 2309.69213867188, 
    2309.69213867188, 1210.18420410156, 1438.15112304688, 3121.66577148438, 
    3291.59228515625, 3225, 3225, 3550, 3550, 4150, 4150, 4758.9638671875, 
    4758.9638671875, 4694.77685546875, 4384.07421875, 4234.69287109375, 
    4130.41455078125, 4352.24853515625, 4351.2958984375, 4208.11767578125, 
    4326.75439453125, 4260.1845703125, 4137.849609375, 4129.91064453125, 
    3992.22680664062, 3835.96508789062, 3722.62670898438, 3727.2236328125, 
    3425.12133789062, 3236.76147460938, 3221.51342773438, 3115.0966796875, 
    2957.37133789062, 2704.35327148438, 2200.34936523438, 2082.275390625, 
    2211.82006835938, 2385.45336914062, 2524.81079101562, 2620.08422851562, 
    2687.52856445312, 2701.68872070312, 2835.77197265625, 2768.53833007812, 
    2378.57397460938, 2409.95825195312, 3170, 3170, 3178.04028320312, 
    3289.48315429688, 3289.48315429688, 3351.72583007812, 3614.56201171875, 
    4043.46752929688, 3913.7236328125, 3786.14697265625, 3398.2001953125, 
    3312.47241210938, 3312.47241210938, 3139.02783203125, 3264.02490234375, 
    3010, 3016.24291992188, 3376.4033203125, 3372.24438476562, 
    3323.48779296875, 4557.74462890625, 4695.9453125, 4850.4296875, 
    5445.19482421875, 5258.9287109375, 5352.314453125, 5390.77099609375, 
    5184.9384765625, 4590.5166015625, 4639.3134765625, 4406.27099609375, 
    3839.0185546875, 2804.73046875, 2478.65795898438, 2762.44287109375, 
    2997.4306640625, 2916.0771484375, 2440, 2440, 3070.27905273438, 4155, 
    4155, 4155, 4155, 4185, 4185, 4088.33911132812, 4560.13720703125, 
    4528.40283203125, 4365.5029296875, 4403.43359375, 4703.0634765625, 
    5059.9169921875, 4826.43603515625, 4742.466796875, 4638.85400390625, 
    4599.64404296875, 4368.72314453125, 4606.6025390625, 4543.177734375, 
    4400.93017578125, 4225.2744140625, 4045.58276367188, 3504.50439453125, 
    1880.51611328125, 1203.83923339844, 1161.10522460938, 1254.36962890625, 
    1106.42602539062, 1413.08569335938, 1535.29650878906, 1998.08666992188, 
    3445.13403320312,
  3676.73095703125, 3566.916015625, 3989.00317382812, 4350.5146484375, 
    4375.63330078125, 4375.63330078125, 4340.4169921875, 4367.708984375, 
    4367.708984375, 4265.40966796875, 4147.380859375, 4224.48046875, 
    4135.064453125, 4079.38330078125, 3967.77001953125, 3823.05908203125, 
    3874.4638671875, 3838.34545898438, 3873.95874023438, 3704.53149414062, 
    3675.48657226562, 3593.4541015625, 3617.73681640625, 3533.939453125, 
    3452.91479492188, 3656.19604492188, 3655.16625976562, 3655.16625976562, 
    3613.9716796875, 3531.96899414062, 3470.22900390625, 3569.27319335938, 
    3671.31396484375, 3640.9091796875, 3698.98413085938, 3698.98413085938, 
    3876.56030273438, 3873.34375, 4065.89147763595, 4247.28662109375, 
    4379.8564453125, 4351.0283203125, 4351.0283203125, 4342.7470703125, 
    4582.12548828125, 4528.22119140625, 4377.60888671875, 4035.19213867188, 
    3897.4619140625, 3843.82495117188, 3844.02221679688, 3673.3603515625, 
    3601.57885742188, 3432.73559570312, 3459.64379882812, 3423.43041992188, 
    3174.00073242188, 3124.64721679688, 2788.71118164062, 2730.61962890625, 
    2884.0859375, 3079.66723632812, 3333.748046875, 3333.748046875, 
    3257.77661132812, 3292.95141601562, 4050, 4050, 4050, 4050, 4050, 4050, 
    4091.72143554688, 4247.7265625, 4395.96875, 4288.54931640625, 
    4288.54931640625, 4242.96337890625, 4239.23486328125, 3898.25610351562, 
    1971.4453125, 3446.36450195312, 3857.23413085938, 3857.23413085938, 
    3606.22607421875, 1281.94848632812, 1118.384765625, 963.555786132812, 
    425.785466617812, 150, 346.236572265625, 346.236572265625, 
    343.311187744141, 604.643127441406, 3138.10595703125, 4577.56201171875, 
    4978.59521484375, 4998.54150390625, 5000.541015625, 5056.93017578125, 
    5064.84912109375, 5279.45947265625, 5346.52001953125, 5479.12158203125, 
    5500, 5500, 5500, 5500, 5500, 5409.93359375, 5265.109375, 5272.484375, 
    5125.15087890625, 5089.8017578125, 4919.94775390625, 4851.24560546875, 
    4764.30712890625, 4725.103515625, 4536.8798828125, 4520.85791015625, 
    4333.15771484375, 4229.83349609375, 4309.65283203125, 4320, 
    4309.45654296875, 4309.45654296875, 4166.54833984375, 4310.76611328125, 
    4379.27734375, 4379.27734375, 4311.33154296875, 4394.83447265625, 
    4114.6962890625, 3973.06713867188, 3866.70336914062, 3927.43017578125, 
    3721.27612304688, 2704.5263671875, 3078.58740234375, 3577.74267578125, 
    3577.74267578125, 3459.88403320312, 4209.17919921875, 4209.3935546875, 
    4404.41552734375, 4335.60546875, 4342.38916015625, 4361.02978515625, 
    4042.04907226562, 4002.83129882812, 4032.43115234375, 4032.43115234375, 
    3864.76123046875, 3795.775390625, 3578.259765625, 3489.67358398438, 
    3350.12255859375, 3275.24340820312, 3107.22436523438, 2816.05419921875, 
    2687.4423828125, 2604.31176757812, 2722.02465820312, 3025.84033203125, 
    3285.63793945312, 3442.96655273438, 3539.63647460938, 3648.80908203125, 
    3667.22338867188, 3721.27612304688, 3810.62548828125, 3818.84716796875, 
    3927.94091796875, 3986.35766601562, 4135.05859375, 4232.8173828125, 
    4165.17529296875, 4256.60400390625, 4360.6328125, 4360.6328125, 
    4380.14208984375, 4545.89990234375, 4647.9833984375, 4605.978515625, 
    4678.474609375, 4671.84375, 4880.27978515625, 4883.4765625, 
    4921.7763671875, 4912.27294921875, 4912.54833984375, 4878.35888671875, 
    4842.7978515625, 4839.431640625, 4851.26513671875, 4719.94091796875, 
    4558.95361328125, 4462.78466796875, 4371.0546875, 4226.890625, 
    4075.66870117188, 3917.20629882812, 4000.76904296875, 3969.63549804688, 
    561.327819824219, 0, -0, -0, -0, -0, -0, 40, 90, 110, 130, 150, 
    257.514770507812, 311.124694824219, 313.010345458984, 170, 60, 140, 
    426.629821777344, 1297.03967285156, 1592.55358886719, 1974.64294433594, 
    1974.64294433594, 2072.27514648438, 2274.41650390625, 2337.615234375, 
    2417.87719726562, 3252.77490234375, 3252.77490234375, 2651.83740234375, 
    2651.83740234375, 2651.83740234375, 2232.54907226562, 1814.62548828125, 
    2948.19848632812, 3699.1318359375, 3699.1318359375, 3479.17333984375, 
    2620.9609375, 3010.4765625, 3835.29833984375, 3751.82885742188, 3050, 
    3050, 3245.55102539062, 3245.55102539062, 4150, 4120.5537109375, 
    4685.11865234375, 4435.2275390625, 4150, 3041.84448242188, 
    4208.79541015625, 4237.89501953125, 4274.47509765625, 4274.47509765625, 
    4263.81103515625, 4278.57080078125, 4225.7939453125, 4162.154296875, 
    4039.23950195312, 3957.28491210938, 3866.95556640625, 3648.02392578125, 
    3677.96435546875, 3416.86938476562, 3042.05346679688, 2814.56323242188, 
    2708.369140625, 2580.9716796875, 2667.32568359375, 2432.04516601562, 
    2449.58129882812, 2446.88354492188, 2450.73828125, 2573.59252929688, 
    2745.00170898438, 2615.62475585938, 2565.04272460938, 2768.53833007812, 
    3367.31860351562, 3656.78173828125, 3538.16528320312, 3575.708984375, 
    3520.59887695312, 3287.7431640625, 2955.57983398438, 2863.2880859375, 
    3180.20043945312, 3180.20043945312, 2733.42114257812, 2924.8916015625, 
    3007.99780273438, 3010, 3010, 3010, 3010, 3010, 2959.30737304688, 
    2959.30737304688, 3557.42431640625, 3557.42431640625, 3459.97631835938, 
    3249.29833984375, 4529.8779296875, 4844.6728515625, 5131.455078125, 5500, 
    5384.47216796875, 5254.875, 5175.1904296875, 4500.4619140625, 
    4454.53564453125, 4356.2822265625, 4070.28271484375, 3370.859375, 
    2547.62768554688, 1920, 2281.29248046875, 2281.29248046875, 2100, 
    3175.70678710938, 3079.91796875, 4155, 4155, 4155, 4185, 4503.5732421875, 
    4503.5732421875, 4085.39453125, 4225, 4312.60498046875, 4365.5029296875, 
    4664.6982421875, 4703.0634765625, 4926.72998046875, 4896.32958984375, 
    4567.63720703125, 4584.01708984375, 4501.22607421875, 4368.72314453125, 
    4368.72314453125, 4334.01708984375, 4069.41162109375, 3878.3525390625, 
    3802.97607421875, 3156.29467773438, 1579.47485351562, 409.609832763672, 
    220, 230, 539.122497558594, 664.960632324219, 1172.60766601562, 
    2345.15112304688, 3639.203125,
  3722.896484375, 3877.25537109375, 4031.6474609375, 4249.39892578125, 
    4311.52392578125, 4257.1494140625, 4206.85986328125, 4302.59765625, 
    4285.5498046875, 4150.97314453125, 4157.15576171875, 4188.888671875, 
    4023.6318359375, 4040.17358398438, 3938.07836914062, 3864.74658203125, 
    3852.4697265625, 3750.40649414062, 3725.46484375, 3694.07934570312, 
    3638.84301757812, 3587.0966796875, 3579.57861328125, 3515.85498046875, 
    3473.76684570312, 3460.0224609375, 3597.3466796875, 3586.15502929688, 
    3535.4736328125, 3387.2978515625, 3479.76635742188, 3569.27319335938, 
    3591.2353515625, 3542.2177734375, 3603.12329101562, 3700.20874023438, 
    3698.98413085938, 3659.27392578125, 3675.68432617188, 3866.8466796875, 
    4114.7880859375, 4249.97900390625, 4398.55029296875, 4205.07275390625, 
    4045, 4194.43115234375, 4139.7607421875, 3829.7568359375, 
    3604.94677734375, 3625.98364257812, 3603.427734375, 3423.978515625, 
    3387.2978515625, 3371.07568359375, 3265.7041015625, 3258.38891601562, 
    3178.39990234375, 3032.88208007812, 2690.30834960938, 2737.4228515625, 
    3492.71655273438, 3625.22729492188, 3653.26196289062, 4155, 4155, 4155, 
    4080.99853515625, 4067.38598632812, 4226.80078125, 4050, 4050, 
    4151.8310546875, 4289.833984375, 4351.53662109375, 4380.48974609375, 
    4380.48974609375, 4380.48974609375, 4335.0244140625, 4310.86376953125, 
    3898.25610351562, 3499.73291015625, 2441.18896484375, 3488.57592773438, 
    3606.22607421875, 3606.22607421875, 1159.69897460938, 692.589599609375, 
    632.42236328125, 470.114532470703, 470.114532470703, 484.749450683594, 
    484.749450683594, 457.117004394531, 634.507385253906, 814.675842285156, 
    2665.87890625, 4732.6494140625, 4998.4931640625, 4879.2900390625, 
    4936.89404296875, 4874.212890625, 4975.6943359375, 5036.66552734375, 
    5146.97119140625, 5403.6630859375, 5277.859375, 5500, 5317.91064453125, 
    5096.90234375, 5096.90234375, 5022.75390625, 5125.15087890625, 
    5125.15087890625, 5089.8017578125, 4948.5595703125, 4888.97412109375, 
    4803.9287109375, 4927.49658203125, 4722.02587890625, 4563.345703125, 
    4605.4443359375, 4367.62109375, 4539.63623046875, 4539.63623046875, 
    4400.9140625, 4309.45654296875, 4460.33447265625, 4644.44775390625, 
    4601.474609375, 4437.37646484375, 4311.33154296875, 4280.19189453125, 
    4264.3466796875, 4037.55786132812, 3925.97924804688, 4027.3623046875, 
    4027.3623046875, 3981.59326171875, 3582.07202148438, 4123.83056640625, 
    4403.859375, 4271.04443359375, 4209.17919921875, 4408.79443359375, 
    4209.3935546875, 4383.228515625, 4363.3408203125, 4539.67236328125, 
    4419.18185522252, 4206.9248046875, 4166.81689453125, 4032.43115234375, 
    3960.96459960938, 3777.275390625, 3647.90405273438, 3529.84619140625, 
    3544.91748046875, 3532.62036132812, 3326.11669921875, 3169.58862304688, 
    2997.38452148438, 2847.97924804688, 2730.65625, 3048.06176757812, 
    3199.06713867188, 3387.2978515625, 3484.66455078125, 3534.94921875, 
    3667.22338867188, 3745.69750976562, 3739.44921875, 3818.9384765625, 
    3823.41674804688, 3907.67041015625, 4050.27661132812, 4050.27661132812, 
    4106.29296875, 4200.46826171875, 4360.6328125, 4360.6328125, 
    4399.87158203125, 4535.962890625, 4627.33349609375, 4628.126953125, 
    4671.84375, 4892.79345703125, 4901.31689453125, 4842.1796875, 
    4819.95947265625, 4792.42236328125, 4728.06689453125, 4733.92724609375, 
    4655.13916015625, 4588.17041015625, 4437.4755859375, 4342.71875, 
    4238.95947265625, 4379.740234375, 4287.283203125, 4031.93505859375, 
    3888.64697265625, 3885.20361328125, 3937.72900390625, 3561.70190429688, 
    550, 0, -0, -0, -0, -0, -0, 50, 90, 120, 130, 150, 180, 180, 120, 0, -0, 
    -0, 120, 603.885681152344, 1145.75048828125, 1551.9609375, 
    1862.40393066406, 2072.27514648438, 2274.41650390625, 2337.615234375, 
    2417.87719726562, 2450.11938476562, 2621.6728515625, 2735.7724609375, 
    2651.83740234375, 2683.20239257812, 2232.54907226562, 1814.62548828125, 
    2948.19848632812, 3699.1318359375, 3735.46313476562, 4003.00439453125, 
    4405.26416015625, 4405.26416015625, 3751.82885742188, 3751.82885742188, 
    3050, 3040.17041015625, 3536.80590820312, 4150, 4150, 4407.2119140625, 
    4211.876953125, 3250, 3250, 4282.08251953125, 4498.17041015625, 
    4607.6220703125, 4496.1904296875, 4301.33642578125, 4398.42919921875, 
    4402.43798828125, 4313.859375, 4315.81640625, 4039.23950195312, 
    3461.13671875, 3778.21923828125, 3789.17309570312, 3694.07543945312, 
    3625.76513671875, 3029.9462890625, 2625.33911132812, 2558.54907226562, 
    2227.36328125, 2066.77514648438, 2358.93823242188, 2664.26782226562, 
    2819.45947265625, 2891.52587890625, 2683.34545898438, 2155.81225585938, 
    2867.27124023438, 2867.27124023438, 2767.82421875, 3367.31860351562, 
    3538.16528320312, 3807.87744140625, 3906.59936523438, 3943.77124023438, 
    4036.6767578125, 3763.52368164062, 3306.68579101562, 2475.12963867188, 
    2970.73193359375, 3367.68627929688, 3166.57495117188, 3333.03369140625, 
    3431.01123046875, 3402.91333007812, 3595.6416015625, 3595.6416015625, 
    3688.69067382812, 3688.69067382812, 4017.80810546875, 3917.03149414062, 
    3971.39599609375, 3971.39599609375, 3835.46508789062, 4294.7548828125, 
    4346.47802734375, 4850, 5021.998046875, 5021.998046875, 4951.232421875, 
    4945.39453125, 4737.873046875, 4636.6162109375, 4407.4169921875, 
    4082.48388671875, 3464.1005859375, 3216.71435546875, 3150, 3150, 3150, 
    3167.55444335938, 3648.763671875, 3800.68188476562, 4156.03369140625, 
    4507.37451171875, 4614.771484375, 4379.443359375, 4531.90576171875, 
    4529.29541015625, 4463.18994140625, 4225, 4225, 4348.41796875, 
    4597.91650390625, 4703.0634765625, 4734.625, 4545.34033203125, 4545, 
    4552.1484375, 4385.66845703125, 4190.48828125, 3622.20629882812, 
    2966.10034179688, 2284.19116210938, 2284.19116210938, 2169.06079101562, 
    633.14013671875, 640, 640, 640, 425.785466617812, 556.317199707031, 
    1960.2216796875, 3204.8642578125, 3555.77221679688, 3640,
  3879.56787109375, 3967.49072265625, 4031.6474609375, 4193.57666015625, 
    4218.9716796875, 4188.99072265625, 4220.62841796875, 4137.1552734375, 
    4065.89147763595, 4102.73779296875, 4042.5390625, 3966.29931640625, 
    3837.91772460938, 3775.60620117188, 3666.10083007812, 3608.8544921875, 
    3628.00073242188, 3672.35302734375, 3570.892578125, 3518.55126953125, 
    3618.45581054688, 3641.83666992188, 3524.33374023438, 3264.7451171875, 
    3294.97583007812, 3338.26782226562, 3344.32373046875, 3237.09057617188, 
    3227.97827148438, 3170.30908203125, 3300.73364257812, 3300.73364257812, 
    3291.62280273438, 3264.9384765625, 3426.25756835938, 3639.14306640625, 
    3639.14306640625, 3552.14013671875, 3492.74340820312, 3442.21508789062, 
    3681.30102539062, 3674.59643554688, 3706.10424804688, 4051.52368164062, 
    4045, 4072.41088867188, 4261.79150390625, 3444.45654296875, 
    3452.4091796875, 3371.33959960938, 3283.12890625, 3222.94873046875, 
    3202.49291992188, 2959.13110351562, 2977.64770507812, 2949.6064453125, 
    3029.56030273438, 3030, 3030, 3193.06201171875, 3642.84375, 3642.84375, 
    4155, 4155, 4155, 4155, 4155, 4231.71240234375, 4380.49267578125, 4050, 
    4050, 4257.83056640625, 4354.1552734375, 4351.53662109375, 
    4419.64404296875, 4598.22412109375, 4481.61572265625, 4422.505859375, 
    4393.341796875, 4250.01904296875, 4080.09619140625, 3919.78784179688, 
    1766, 1684.53723144531, 2399.29858398438, 2399.29858398438, 80, 
    309.836761474609, 556.824462890625, 567.390258789062, 568.238464355469, 
    484.749450683594, 457.117004394531, 605.291259765625, 814.675842285156, 
    1600.32397460938, 2953.78295898438, 3790.10620117188, 4325.21728515625, 
    4383.58154296875, 4383.58154296875, 4253.021484375, 3468.9501953125, 
    4400, 5011.92333984375, 5332.61962890625, 5390.14599609375, 
    5143.41858983545, 5073.08740234375, 5112.55029296875, 5074.654296875, 
    5117.50732421875, 5057.322265625, 5114.8505859375, 5114.8505859375, 
    5114.07568359375, 5103.806640625, 4929.771484375, 4804.7607421875, 
    4703.55908203125, 4991.72802734375, 5085.966796875, 4970.1455078125, 
    5005.27734375, 4880.7490234375, 4583.150390625, 4745.6337890625, 
    4726.71435546875, 4684.474609375, 4548.552734375, 4311.33154296875, 
    4312.74365234375, 4320, 4327.2197265625, 4327.2197265625, 
    4135.66650390625, 4158.96826171875, 4763.478515625, 4643.080078125, 
    4506.75, 4065.89147763595, 4272.00537109375, 4408.55712890625, 
    4408.55712890625, 4599.6640625, 4555.04638671875, 4642.5517578125, 
    4598.7822265625, 4532.0517578125, 4327.07666015625, 4110.22412109375, 
    4007.03198242188, 3960.96459960938, 3879.7099609375, 3687.76513671875, 
    3631.6318359375, 3564.69653320312, 3513.15649414062, 3326.11669921875, 
    3259.35107421875, 3122.17724609375, 2873.51538085938, 2730.65625, 
    2832.5830078125, 2918.78759765625, 3115.568359375, 3258.42016601562, 
    3456.79345703125, 3574.61938476562, 3611.82958984375, 3492.2119140625, 
    3681.29736328125, 3786.25463867188, 3850.26147460938, 4013.8876953125, 
    3998.03100585938, 4145.9970703125, 4216.73193359375, 4214.76513671875, 
    4345.869140625, 4271.26318359375, 4262.9541015625, 4190.28466796875, 
    4505.65478515625, 4647.69970703125, 4855.0244140625, 4995.23095703125, 
    4867.1669921875, 4841.5703125, 4764.0947265625, 4752.78515625, 
    4634.86181640625, 4586.52685546875, 4485.16162109375, 4438.4345703125, 
    4397.41259765625, 4362.96630859375, 4272.99853515625, 4194.89501953125, 
    4018.7822265625, 3906.84350585938, 3870.984375, 3957.16455078125, 
    1839.66296386719, 0, -0, -0, -0, -0, -0, -0, 50, 60, 120, 120, 150, 150, 
    150, 150, 150, 160, 160, 253.361404418945, 495.553629324057, 
    942.839303029559, 1381.59167480469, 1807.28454589844, 2046.53198242188, 
    2149.74072265625, 2316.02001953125, 2720.21655273438, 2721.18334960938, 
    2721.18334960938, 2156.35424804688, 1827.87780761719, 1506.20056152344, 
    1423.97717285156, 1452.52124023438, 1768.38269042969, 2506.71533203125, 
    4021.63989257812, 4877.9462890625, 5025.14208984375, 4605.7119140625, 
    3619.51489257812, 4710.07275390625, 4586.38623046875, 4631.49755859375, 
    4710.4765625, 4843.67041015625, 4914.3046875, 4211.876953125, 
    4211.876953125, 3253.5576171875, 3807.650390625, 4542.828125, 
    4470.61474609375, 4452.4404296875, 4454.83447265625, 4301.33642578125, 
    4361.64306640625, 4388.6171875, 4277.10498046875, 4148.76708984375, 
    3959.01684570312, 3721.27612304688, 3730.81420898438, 3875.8837890625, 
    3441.44384765625, 3387.2978515625, 3029.9462890625, 2655.23876953125, 
    2386.10522460938, 2483.43676757812, 2599.07006835938, 2636.95849609375, 
    2743.7265625, 2813.01684570312, 2894.19189453125, 2584.01708984375, 
    3327.42993164062, 3396.29028320312, 3423.69091796875, 2275.8828125, 
    2926.66723632812, 2926.66723632812, 3744.11791992188, 4008.06713867188, 
    4213.33203125, 4238.3037109375, 3871.04174804688, 3490.38208007812, 
    3490.38208007812, 3069.51513671875, 3620.57202148438, 3875.92260742188, 
    3974.45776367188, 4027.28076171875, 4027.28076171875, 3857.33471679688, 
    4143.97607421875, 4190.068359375, 4190.068359375, 4174.623046875, 
    4174.623046875, 4175, 4175, 4260, 4260, 4260, 4260, 4831.36083984375, 
    4931.2353515625, 4931.2353515625, 4931.2353515625, 4737.873046875, 
    4636.6162109375, 4347.033203125, 4201.9931640625, 3966.11303710938, 
    3807.23095703125, 3810, 3944.486328125, 4136.2099609375, 4066.8525390625, 
    4093.22290039062, 4373.69384765625, 4246.4189453125, 4584.654296875, 
    4534.76806640625, 4379.443359375, 4449.24755859375, 4666.3935546875, 
    4543.1484375, 4271.06689453125, 4283.83984375, 4152.7119140625, 
    4451.4130859375, 4629.1220703125, 4629.1220703125, 4545, 4545, 
    4598.49609375, 4123.93798828125, 2449.13256835938, 2467.72265625, 
    2487.236328125, 1753.32263183594, 1361.45544433594, 468.865447998047, 
    640.254150390625, 640, 640, 640, 838.071899414062, 1631.00854492188, 
    2899.2060546875, 3467.0625, 3526.94165039062, 3637.60083007812,
  3786.01904296875, 3724.49853515625, 3941.09008789062, 4099.5029296875, 
    4125.33544921875, 4185.267578125, 4047.09326171875, 4048.01025390625, 
    4048.01025390625, 3982.81127929688, 3965.37036132812, 3792.43090820312, 
    3805.56616210938, 3622.70581054688, 3552.9033203125, 3493.48559570312, 
    3260, 3260, 3260, 3268.51782226562, 3358.58740234375, 3314.076171875, 
    3312.29077148438, 3181.11791992188, 3161.662109375, 3115.27319335938, 
    3019.66967773438, 3267.79345703125, 3261.76513671875, 3193.96435546875, 
    3133.22705078125, 3239.88208007812, 3440.11840820312, 3547.349609375, 
    3374.92797851562, 3598.53735351562, 3569.283203125, 3590.9375, 
    3548.91821289062, 3605.10278320312, 3984.13134765625, 3814.70874023438, 
    3527.38549804688, 4045, 4045, 4045, 4045, 3824.93530273438, 
    3733.14916992188, 3676.7861328125, 3684.59252929688, 3558.28051757812, 
    3527.63452148438, 3404.94970703125, 3352.60864257812, 3438.0673828125, 
    3464.5859375, 3253.53393554688, 3130.52490234375, 3149.10693359375, 
    3642.84375, 4155, 4155, 4155, 4155, 4387.5537109375, 4108.6767578125, 
    4325.986328125, 4196.96142578125, 3197.13110351562, 2570.51000976562, 
    4165, 4369.197265625, 4346.54052734375, 4670.037109375, 4586.484375, 
    4556.06005859375, 4747.6103515625, 4747.6103515625, 4546.8212890625, 
    4346.130859375, 4186.57470703125, 3701.58227539062, 3701.58227539062, 
    2399.29858398438, 2399.29858398438, 326.990295410156, 309.836761474609, 
    664.199645996094, 665.210815429688, 563.388732910156, 333.346130371094, 
    430.907928466797, 495.573974609375, 516.286254882812, 1050, 1050, 
    955.042541503906, 879.3212890625, 1742.07043457031, 2994.55029296875, 
    3436.56494140625, 3436.56494140625, 4400, 5072.734375, 5335.1875, 
    5370.98046875, 5326.78466796875, 5240.2890625, 5183.3603515625, 
    5242.099609375, 5322.57958984375, 5251.56103515625, 5145.3583984375, 
    5237.0400390625, 5114.07568359375, 5108.66357421875, 4945.716796875, 
    4878.60205078125, 5027.07373046875, 4991.72802734375, 5072.375, 
    5032.16796875, 5020.56103515625, 5103.57373046875, 4749.52734375, 
    4749.52734375, 4750.59619140625, 4498.20556640625, 4483.91015625, 
    4191.25390625, 4308.8603515625, 4656.11474609375, 4575.81640625, 
    4515.5361328125, 4566.94775390625, 4531.541015625, 4515.47509765625, 
    4662.19921875, 4504.35546875, 4387.41455078125, 4750.23046875, 
    4426.8408203125, 4491.16650390625, 4680.24267578125, 4739.38330078125, 
    4739.38330078125, 4513.44580078125, 4532.19482421875, 4336.16845703125, 
    4110.67236328125, 3942.18310546875, 3975.97778320312, 3913.25512695312, 
    3915.73901367188, 3823.99731445312, 3652.28100585938, 3480.18286132812, 
    3226.26513671875, 3216.29296875, 3076.18505859375, 2846.716796875, 
    2679.25634765625, 2868.60620117188, 2904.82592773438, 2904.82592773438, 
    2658.90698242188, 2942.55541992188, 3110.40551757812, 3256.68872070312, 
    3397.28198242188, 3593.14990234375, 3771.73120117188, 3821.9599609375, 
    3869.2998046875, 4035.23364257812, 4019.28955078125, 4150.8125, 
    4242.0556640625, 4324.11962890625, 4308.95068359375, 4329.90576171875, 
    4321.2890625, 4517.24853515625, 4631.47900390625, 4779.07571895829, 
    4896.4248046875, 4736.7314453125, 4706.2021484375, 4645.66552734375, 
    4663.052734375, 4604.79150390625, 4490.23974609375, 4471.89306640625, 
    4397.47802734375, 4362.96630859375, 4362.96630859375, 4173.8818359375, 
    4097.7255859375, 3987.45727539062, 3836.78735351562, 3891.73217773438, 
    3973.25415039062, 1935.05359591651, 0, -0, -0, -0, -0, -0, -0, -0, 40, 
    110, 120, 140, 150, 150, 160, 200, 345.196807861328, 348.018035888672, 
    348.018035888672, 646.283386230469, 980.161560058594, 1302.18920898438, 
    1886.43371582031, 2476.30834960938, 3311.58764648438, 3621.341796875, 
    4663.01171875, 4610.892578125, 4641.91259765625, 4491.087890625, 
    4663.62939453125, 4663.62939453125, 4136.80517578125, 3750.373046875, 
    3430.349609375, 3355.9052734375, 4021.63989257812, 4779.07571895829, 
    5085.05810546875, 4960.2783203125, 5077.55322265625, 5111.6015625, 4965, 
    4754.4912109375, 4710.4765625, 5007.859375, 4930.41552734375, 4150, 
    3958.48095703125, 4586.6826171875, 4606.03857421875, 4650.9326171875, 
    4451.79443359375, 4310.5595703125, 4150, 4077.39086914062, 
    4260.9267578125, 4204.982421875, 4183.40966796875, 4100.9931640625, 
    3937.1259765625, 3721.27612304688, 3591.40869140625, 3524.9814453125, 
    3354.67431640625, 3241.51977539062, 2981.94921875, 2655.23876953125, 
    2976.5078125, 2939.494140625, 3214.74096679688, 3430.46630859375, 
    3520.81958007812, 3368.05981445312, 3406.98559570312, 3578.25805664062, 
    3727.89086914062, 3844.58935546875, 3662.24438476562, 3668.33935546875, 
    3402.09155273438, 3229.06323242188, 2758.41088867188, 1960.03881835938, 
    4089.01123046875, 4191.43310546875, 3842.71313476562, 3924.03637695312, 
    3822.90625, 4046.72607421875, 4046.72607421875, 4328.27880859375, 
    4328.27880859375, 4328.27880859375, 4232.3427734375, 4238.560546875, 
    4288.29541015625, 4288.29541015625, 4252.37646484375, 4490.00634765625, 
    4757.484375, 4747.6533203125, 4747.6533203125, 4720.07666015625, 
    4450.6435546875, 4260, 4260, 4175, 4343.5390625, 4700.46240234375, 
    4504.2919921875, 4506.80224609375, 4290.046875, 4323.8359375, 
    4323.8359375, 4406.4423828125, 4246.08837890625, 4198.80078125, 
    4047.02563476562, 4239.564453125, 4372.25927734375, 4306.04931640625, 
    4346.38916015625, 4246.4189453125, 4162.38623046875, 4238.1142578125, 
    4263.4560546875, 4292.3486328125, 4312.04345703125, 4338.244140625, 
    4294.021484375, 4255.53076171875, 4317.0986328125, 4460.041015625, 
    4504.3046875, 4599.01904296875, 4524.06005859375, 3485.41625976562, 
    3225.66748046875, 1644.84631347656, 1634.64953613281, 1634.64953613281, 
    1579.4462890625, 387.202423095703, 90, -0, 90, 580.953491210938, 
    1284.98950195312, 2175.3212890625, 2568.25, 2902.87548828125, 
    3131.65454101562, 3415.3818359375, 3512.26928710938, 3640.58203125,
  3581.18530273438, 3520.90356445312, 3668.46215820312, 3828.24780273438, 
    3980.35180664062, 4019.01147460938, 4005.94409179688, 3792.67456054688, 
    3893.671875, 3864.21997070312, 3776.46166992188, 3849.02075195312, 
    3697.44677734375, 3326.21069335938, 3326.21069335938, 3314.34204101562, 
    3214.525390625, 3009.876953125, 3050, 3067.197265625, 3125.98291015625, 
    3088.03833007812, 3164.75415039062, 3150.45971679688, 3001.962890625, 
    3126.05590820312, 3088.01904296875, 2954.40551757812, 3188.87890625, 
    3519.0771484375, 3557.37646484375, 3509.22583007812, 3581.65209960938, 
    3641.57153320312, 3641.57153320312, 3689.97021484375, 3561.48510742188, 
    3826.37158203125, 3840.06591796875, 3833.53247070312, 3892.59594726562, 
    4046.82543945312, 3911.81640625, 4045, 4045, 4045, 4045, 
    3889.60791015625, 3939.19458007812, 3958.728515625, 3862.80541992188, 
    3810.11547851562, 3837.81787109375, 3693.3857421875, 3611.107421875, 
    3652.49462890625, 3652.49462890625, 3598.42236328125, 3514.40576171875, 
    3651.92236328125, 4278.9130859375, 4133.6259765625, 4158.10888671875, 
    4155, 4155, 4155, 2845.34741210938, 2912.11474609375, 2655.91235351562, 
    1854.48352050781, 1898.70251464844, 4178.6376953125, 4581.20751953125, 
    4581.20751953125, 4642.3671875, 4692.94970703125, 4692.94970703125, 
    4747.6103515625, 4747.6103515625, 4700.10986328125, 4503.30078125, 
    4400.96435546875, 3701.58227539062, 3880.46337890625, 3880.46337890625, 
    2834.876953125, 326.990295410156, 160, 657.746826171875, 
    657.746826171875, 908.875671386719, 908.875671386719, 881.102172851562, 
    867.3779296875, 920.848876953125, 1050, 1050, 955.042541503906, 
    792.583801269531, 657.790954589844, 912.915649414062, 3436.56494140625, 
    4660.0029296875, 4927.97021484375, 5091.55419921875, 5256.55517578125, 
    5390.9482421875, 5373.494140625, 5313.60546875, 5271.2548828125, 
    5307.4404296875, 5281.849609375, 5186.376953125, 5192.005859375, 
    5172.439453125, 5029.8994140625, 4880.5087890625, 4821.86474609375, 
    5038.189453125, 5045.2509765625, 4981.91748046875, 4978.494140625, 
    4921.29443359375, 4839.3076171875, 4790.357421875, 4749.52734375, 
    4753.615234375, 4678.708984375, 4647.79345703125, 4587.1923828125, 
    4682.0517578125, 4308.8603515625, 4534.5068359375, 4429.20703125, 
    4673.01416015625, 4691.21484375, 4529.00244140625, 4731.60400390625, 
    4742.51318359375, 4742.51318359375, 4721.7216796875, 4677.5419921875, 
    4674.80615234375, 4678.078125, 4758.56884765625, 4752.07275390625, 
    4739.38330078125, 4609.28662109375, 4475.87548828125, 4419.18185522252, 
    4419.18185522252, 4204.38427734375, 4102.57275390625, 3913.25512695312, 
    3777.1904296875, 3748.27905273438, 3767.3037109375, 3615.86352539062, 
    3709.26489257812, 3624.14868164062, 3472.00805664062, 3168.57861328125, 
    2985.5810546875, 3053.53247070312, 3012.84033203125, 2767.7705078125, 
    2603.96362304688, 2851.11108398438, 3033.01708984375, 3246.2822265625, 
    3364.80590820312, 3600.14453125, 3790.09521484375, 3870.283203125, 
    3960.41284179688, 4004.68139648438, 4136.3427734375, 4242.26708984375, 
    4340.44287109375, 4272.232421875, 4308.95068359375, 4363.63916015625, 
    4332.24462890625, 4626.35498046875, 4686.5244140625, 4678.12548828125, 
    4605.9697265625, 4578.7607421875, 4565.49365234375, 4458.20166015625, 
    4589.66064453125, 4492.919921875, 4473.357421875, 4369.48095703125, 
    4149.10791015625, 4358.19091796875, 4244.91015625, 4144.53271484375, 
    4095.251953125, 3987.45727539062, 4022.29833984375, 3781.1865234375, 
    3925.20434570312, 1935.05359591651, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    40, 100, 120, 130, 150, 160, 355.639770507812, 570.739868164062, 
    1041.32250976562, 1158.96691894531, 1333.61352539062, 2335.20581054688, 
    4420.603515625, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5492.49267578125, 
    5404.3955078125, 5432.44140625, 4965, 4965, 4754.4912109375, 
    4334.16259765625, 4602.14111328125, 4460.41357421875, 4188.9775390625, 
    4651.72412109375, 4541.67138671875, 4438.24658203125, 4335.75830078125, 
    4401.625, 4334.22607421875, 4180.734375, 4065.89147763595, 
    4244.15771484375, 4125.009765625, 3824.92602539062, 3786.27661132812, 
    3615.57543945312, 3621.63623046875, 3338.6865234375, 3023.96704101562, 
    2776.63037109375, 2396.24438476562, 2517.82299804688, 2939.4814453125, 
    3375.33642578125, 3612.59521484375, 3604.9345703125, 3746.529296875, 
    3788.63452148438, 3945.34423828125, 3726.31005859375, 3701.294921875, 
    3756.62573242188, 3722.3818359375, 4009.9716796875, 4009.9716796875, 
    3901.67407226562, 3160.94506835938, 3177.630859375, 2172.45776367188, 
    3306.89819335938, 3289.71166992188, 3954.37744140625, 3791.31665039062, 
    3961.52099609375, 4212.92041015625, 4649.55810546875, 4649.55810546875, 
    4390.87060546875, 4701.08740234375, 4701.08740234375, 4675.0849609375, 
    4538.951171875, 4383.43310546875, 4629.86572265625, 4864.6494140625, 
    4839.27783203125, 5087.22119140625, 5087.22119140625, 4814.46923828125, 
    4814.46923828125, 4319.853515625, 4284.14013671875, 3631.79443359375, 
    3842.4208984375, 4097.74658203125, 4097.74658203125, 4369.22265625, 
    4392.42724609375, 4323.8359375, 4379.1953125, 4212.83154296875, 
    4212.83154296875, 4166.0810546875, 4047.02563476562, 4288.2021484375, 
    4108.89892578125, 4008.60229492188, 4007.50122070312, 3932.13330078125, 
    4044.31982421875, 4137.4365234375, 4065.89147763595, 3960.64819335938, 
    3945.1884765625, 3973.16943359375, 4096.28759765625, 4233.9521484375, 
    4301.166015625, 4397.8125, 4397.8125, 4384.74951171875, 4382.42626953125, 
    3422.99926757812, 2257.271484375, 2329.85278320312, 2329.85278320312, 
    1486.16943359375, 878.186706542969, 253.361404418945, 130, 70, 120, 
    580.953491210938, 1504.55908203125, 2361.3662109375, 2618.30517578125, 
    2957.21118164062, 3103.35717773438, 3271.52075195312, 3352.89965820312, 
    3352.89965820312,
  3426.01782226562, 3387.39111328125, 3525.72924804688, 3668.68896484375, 
    3703.35791015625, 3628.1943359375, 3662.62939453125, 3662.62939453125, 
    3678.7158203125, 3596.48510742188, 3607.0458984375, 3641.50366210938, 
    3696.24755859375, 3389.47729492188, 3326.21069335938, 3082.14868164062, 
    3025, 3025, 2839.14575195312, 2881.6064453125, 2829.994140625, 
    2938.28784179688, 2937.6630859375, 3072.25048828125, 3168.03125, 
    3342.9345703125, 3194.79956054688, 3373.46923828125, 3069.52612304688, 
    3388.49291992188, 3621.68334960938, 3801.4462890625, 3812.91381835938, 
    3929.16040039062, 3923.39697265625, 3984.11767578125, 3837.34204101562, 
    4040.45971679688, 4044.677734375, 3950.97607421875, 4125.50732421875, 
    4246.31103515625, 3911.81640625, 4191.3994140625, 4065.89147763595, 
    4152.04638671875, 4219.72705078125, 4049.77685546875, 4097.32177734375, 
    4197.0244140625, 4096.11474609375, 4122.90087890625, 4086.57958984375, 
    4074.369140625, 4022.35620117188, 4042.94677734375, 3912.04077148438, 
    3863.84545898438, 3815.16625976562, 3934.74584960938, 4153.85888671875, 
    4354.04345703125, 4325.296875, 4155, 4155, 3401.94946289062, 
    2395.35522460938, 1198.99914550781, 1043.17456054688, 2307.02978515625, 
    3204.25048828125, 4341.75341796875, 4581.20751953125, 4753.259765625, 
    4642.3671875, 4692.94970703125, 4692.94970703125, 4672.6025390625, 
    4700.80224609375, 4700.80224609375, 4419.18185522252, 4419.18185522252, 
    4311.9609375, 4304.4765625, 4199.33447265625, 2836.37231445312, 
    595.991271972656, 110, 140, 584.369445800781, 908.875671386719, 
    1264.50268554688, 1390.7138671875, 1397.71350097656, 1249.10925292969, 
    1218.57800292969, 1049.74047851562, 894.533630371094, 595.026733398438, 
    333.937408447266, 994.998657226562, 3167.8935546875, 4660.0029296875, 
    4981.83056640625, 5034.8291015625, 5037.92333984375, 5143.41858983545, 
    5179.72900390625, 5178.845703125, 5228.9384765625, 5146.65673828125, 
    5360.37255859375, 5261.65771484375, 5285.69873046875, 5196.2998046875, 
    5055.197265625, 4836.5712890625, 4865.35693359375, 4713.12158203125, 
    4637.83837890625, 4794.40087890625, 4834.78515625, 4932.15087890625, 
    4931.07666015625, 4817.26220703125, 4756.068359375, 4536.94677734375, 
    4647.79345703125, 4647.79345703125, 4587.1923828125, 4760.38232421875, 
    4767.48681640625, 4751.6357421875, 4751.6357421875, 4434.91943359375, 
    4859.06103515625, 4963.8701171875, 5024.49169921875, 4948.69921875, 
    4884.58642578125, 4979.615234375, 5077.31494140625, 4972.7197265625, 
    5119.42431640625, 4794.048828125, 4768.58837890625, 4696.892578125, 
    4594.5634765625, 4538.923828125, 4468.0380859375, 4419.18185522252, 
    4479.958984375, 4295.68994140625, 4190.16015625, 4177.4423828125, 
    4054.330078125, 3966.92822265625, 3849.24243164062, 3875.36108398438, 
    3770.81787109375, 3659.34057617188, 3490.96923828125, 3263.27172851562, 
    3153.60302734375, 3087.34545898438, 2895.56005859375, 2713.53369140625, 
    2759.90991210938, 2936.92993164062, 3152.69848632812, 3285.8369140625, 
    3499.81372070312, 3621.98071289062, 3721.27612304688, 3920.59619140625, 
    3988.66064453125, 4096.73193359375, 4285.24365234375, 4257.88427734375, 
    4288.888671875, 4374.52783203125, 4141.09716796875, 4391.1630859375, 
    4556.2607421875, 4615.0478515625, 4553.25, 4389.537109375, 
    4389.537109375, 4270.3583984375, 4175, 4172.19091796875, 
    4100.42333984375, 4340.87158203125, 4340.87158203125, 4239.03857421875, 
    3956.96997070312, 3656.42041015625, 3792.27905273438, 3760.34765625, 
    3789.18872070312, 3555.09594726562, 3647.16235351562, 3498.54077148438, 
    3055.7763671875, 485, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 100, 120, 
    130, 130, 355.639770507812, 1041.3955078125, 2505.8837890625, 
    3984.42431640625, 4432.2998046875, 5408.14404296875, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5474.67041015625, 5470.52294921875, 
    5292.49169921875, 5017.1396484375, 4899.00439453125, 4840.3046875, 
    4797.30712890625, 4709.271484375, 4550.32470703125, 4332.96630859375, 
    4406.15771484375, 4403.86572265625, 4230.69482421875, 4255.94384765625, 
    4097.380859375, 3941.53393554688, 3772.69409179688, 3686.19873046875, 
    3571.42431640625, 3308.00952148438, 3065.78548661781, 2939.53881835938, 
    2939.53881835938, 2651.43334960938, 1813.58740234375, 2316.00952148438, 
    3160.72436523438, 3371.7412109375, 3389.74560546875, 3604.9345703125, 
    3845.4794921875, 3971.4033203125, 4000.11596679688, 4026.66748046875, 
    3783.5146484375, 3896.92504882812, 3933.09301757812, 4179.4638671875, 
    4458.6318359375, 4515.154296875, 4290.841796875, 3531.5703125, 
    2172.45776367188, 2887.9091796875, 3250.27880859375, 4297.7236328125, 
    4259.123046875, 4319.2412109375, 4319.2412109375, 4649.55810546875, 
    4711.46142578125, 4534.04052734375, 4701.08740234375, 4936.921875, 
    4936.921875, 5024.06005859375, 4779.07571895829, 4756.013671875, 
    4867.0078125, 5077.59228515625, 5087.22119140625, 5087.22119140625, 
    5422.25390625, 5214.685546875, 4886.4892578125, 4122.65771484375, 
    3436.45336914062, 2432.15698242188, 3251.00659179688, 3251.00659179688, 
    3688.12963867188, 3893.73193359375, 3928.62622070312, 4026.2392578125, 
    4026.2392578125, 3920.87573242188, 3846.02124023438, 3907.11767578125, 
    3262.6103515625, 3654.66821289062, 3503.84399414062, 3241.591796875, 
    3196.60815429688, 3665.70629882812, 3665.70629882812, 3585.39721679688, 
    3639.90014648438, 3692.07983398438, 3692.07983398438, 3875.09106445312, 
    4085.23754882812, 4344.44580078125, 4366.41064453125, 4290.1748046875, 
    4349.005859375, 4349.005859375, 4307.939453125, 3785.85009765625, 
    3666.56298828125, 2871.57958984375, 1571.76000976562, 495.553629324057, 
    331.935119628906, 210, 210, 170, 342.659118652344, 1504.55908203125, 
    2273.09985351562, 2867.07836914062, 3051.58837890625, 3051.80786132812, 
    3304.82080078125, 3233.529296875, 3344.3642578125,
  3437.77685546875, 3411.09326171875, 3555.40307617188, 3576.12329101562, 
    3520.609375, 3626.923828125, 3503.76196289062, 3563.12475585938, 
    3352.8896484375, 3476.96557617188, 3512.8359375, 3434.74096679688, 
    3396.17236328125, 3389.47729492188, 3291.46948242188, 3137.06079101562, 
    3025, 3025, 3102.59399414062, 3131.68188476562, 3008.0546875, 
    3065.78548661781, 3173.43823242188, 3326.67944335938, 3477.53393554688, 
    3575.93408203125, 3611.44702148438, 3598.59692382812, 3569.29663085938, 
    3606.06762695312, 3839.44213867188, 3919.99584960938, 3972.79638671875, 
    3975.2529296875, 3982.611328125, 3988.1357421875, 3969.58447265625, 
    4040.45971679688, 4096.94677734375, 4147.138671875, 4326.462890625, 
    4167.47802734375, 4229.92041015625, 4273.7138671875, 4347.99951171875, 
    4281.2958984375, 4225.9111328125, 4247.953125, 4207.3955078125, 
    4367.31005859375, 4348.62744140625, 4363.619140625, 4332.58837890625, 
    4323.02880859375, 4222.5400390625, 4241.97607421875, 4155, 4155, 4155, 
    4445.26318359375, 4445.6337890625, 4585.10107421875, 4569.1748046875, 
    4155, 3972.31372070312, 3034.75170898438, 2666, 2666, 3535, 4175, 
    4235.212890625, 4563.66162109375, 4526.05078125, 4602.69970703125, 
    4629.83056640625, 4691.48486328125, 4657.75048828125, 4965.12841796875, 
    4880.38232421875, 4990.560546875, 4999.7158203125, 4735.82177734375, 
    4356.86474609375, 4278.3701171875, 4199.33447265625, 2536.45361328125, 
    595.991271972656, 110, 0, -0, 637.883605957031, 1264.50268554688, 
    1420.41052246094, 1420.41052246094, 1308.09875488281, 1401.07348632812, 
    1759.77270507812, 2717.07592773438, 2559.86596679688, 2559.86596679688, 
    2596.80322265625, 3552.53198242188, 4446.7353515625, 4739.400390625, 
    4620.75, 4633.02001953125, 4807.81103515625, 5030.72607421875, 
    5171.892578125, 5255.63330078125, 5404.9912109375, 5410.6787109375, 
    5371.03125, 5403.74951171875, 5268.1669921875, 5212.7822265625, 
    5229.03369140625, 5208.58203125, 4935.3583984375, 4779.07571895829, 
    4715.31640625, 4717.8720703125, 4717.8720703125, 4552.25537109375, 
    4345.37109375, 4692.25146484375, 4619.072265625, 4875.73291015625, 
    4790.2958984375, 4779.07571895829, 4818.375, 4978.28955078125, 
    5064.61962890625, 5037.73828125, 5055.04052734375, 4993.4521484375, 
    5061.58984375, 5061.58984375, 5037.54638671875, 5120.203125, 
    5123.4814453125, 5105.47119140625, 5290.3720703125, 5267.7568359375, 
    4858.92626953125, 4968.970703125, 4862.83447265625, 4690.23583984375, 
    4636.1298828125, 4584.71728515625, 4571.337890625, 4486.80517578125, 
    4456.53759765625, 4311.5546875, 4222.48876953125, 4103.3203125, 
    4033.23681640625, 4033.23681640625, 3968.7802734375, 3781.94580078125, 
    3666.841796875, 3487.23266601562, 3336.74780273438, 3250.93725585938, 
    3099.89038085938, 2947.36743164062, 2713.53369140625, 2859.71118164062, 
    3017.22778320312, 3124.99243164062, 3258.25390625, 3323.08154296875, 
    3323.08154296875, 3454.1640625, 3697.3369140625, 3849.2978515625, 
    3930.13110351562, 4006.05981445312, 4052.12353515625, 4170, 4170, 
    4128.89453125, 4115.78466796875, 4101.7392578125, 4252.68701171875, 
    4312.4775390625, 4170.93310546875, 4150.33251953125, 4146.45166015625, 
    4175, 3958.69970703125, 3721.27612304688, 3981.82666015625, 
    4163.06396484375, 4281.63671875, 3836.91186523438, 3571.13500976562, 
    3656.58959960938, 3286.33715820312, 3555.09594726562, 3555.09594726562, 
    3427.1494140625, 3169.85913085938, 3055.7763671875, 485, -0, -0, -0, -0, 
    -0, -0, -0, -0, 90, 90, 90, 90, 110, 120, 230.335311889648, 
    1127.404296875, 2466.66776221529, 4013.6630859375, 4779.07571895829, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5460.90087890625, 5206.43701171875, 5477.896484375, 5500, 5500, 5500, 
    5329.83349609375, 5500, 5500, 5500, 5500, 5500, 5332.0166015625, 
    5324.8974609375, 5297.994140625, 4910.58837890625, 4905.83447265625, 
    4830.166015625, 4682.54296875, 4767.19970703125, 4464.67431640625, 
    4354.369140625, 4354.369140625, 4152.2724609375, 4141.87646484375, 
    3887.43798828125, 3821.16186523438, 3769.890625, 3463.45288085938, 
    3191.25805664062, 3104.4755859375, 2872.75048828125, 2526.32177734375, 
    2884.56689453125, 2884.56689453125, 2815.05249023438, 3279.5380859375, 
    3279.5380859375, 3122.24462890625, 3681.130859375, 3706.70825195312, 
    3770.0380859375, 3967.04614257812, 4000.11596679688, 4037.6806640625, 
    3914.28930664062, 3896.92504882812, 4126.02294921875, 4605.35205078125, 
    4458.6318359375, 4568.75146484375, 4233.4521484375, 3531.5703125, 
    2524.99047851562, 3707.7900390625, 4679.76318359375, 4741.80615234375, 
    4754.4990234375, 4542.322265625, 4319.2412109375, 4384.2529296875, 
    4556.71875, 4448.69580078125, 4519.26416015625, 4936.921875, 4936.921875, 
    4950.86083984375, 4779.07571895829, 5002.92236328125, 5032.0673828125, 
    5027.7939453125, 5283.99609375, 5500, 5500, 5412.70556640625, 
    5164.775390625, 4851.9345703125, 4482.62109375, 4045.85375976562, 
    3076.39453125, 3331.54931640625, 3069.61767578125, 3018.50024414062, 
    2301.50952148438, 1841.4658203125, 1880.02941894531, 2905.28735351562, 
    2905.28735351562, 1772.26745605469, 2736.03540039062, 2736.03540039062, 
    2069.65185546875, 2106.38037109375, 2747.23364257812, 2747.23364257812, 
    753.735534667969, 570.20361328125, 463.415557861328, 1701.86572265625, 
    3503.11376953125, 3846.82397460938, 4052.80834960938, 4285.7744140625, 
    4454.7578125, 4506.86865234375, 4516.7626953125, 4552.89306640625, 
    4507.1865234375, 4484.8642578125, 4000.6669921875, 3814.85571289062, 
    2805.83837890625, 1416.94213867188, 561.466430664062, 1678.35437011719, 
    2713.46069335938, 2701.0927734375, 2591.26440429688, 3019.50073242188, 
    3463.966796875, 3531.8173828125, 3490.71484375, 3419.46899414062, 
    3402.10107421875, 3513.609375, 3444.53344726562,
  3509.33032226562, 3505.47241210938, 3557.6787109375, 3563.11157226562, 
    3524.50537109375, 3521.06469726562, 3539.48950195312, 3497.95263671875, 
    3352.8896484375, 3310.09375, 3243.1044921875, 3214.05517578125, 
    3115.88647460938, 3228.2412109375, 3134.294921875, 3019.10473632812, 
    3025, 3025, 3348.42993164062, 3389.67309570312, 3410.05126953125, 
    3493.97583007812, 3436.40893554688, 3508.2021484375, 3573.51147460938, 
    3687.087890625, 3814.21606445312, 3947.8173828125, 3779.29345703125, 
    3953.7041015625, 3886.41186523438, 3992.17114257812, 4034.021484375, 
    4023.08520507812, 4120.93994140625, 4105.7958984375, 4164.31103515625, 
    4077.2607421875, 4175.48291015625, 4208.70751953125, 4408.033203125, 
    4242.37939453125, 4435.98583984375, 4462.220703125, 4281.2958984375, 
    4469.76806640625, 4579.38037109375, 4539.8828125, 4419.18185522252, 
    4591.1552734375, 4540.9423828125, 4543.84521484375, 4566.638671875, 
    4484.86865234375, 4419.18185522252, 4396.91162109375, 4321.89208984375, 
    4289.10986328125, 4096.68603515625, 4643.71337890625, 4665.5791015625, 
    4580.5927734375, 4586.75244140625, 4586.75244140625, 3925.75561523438, 
    2666, 2666, 2666, 3535, 4175, 4235.212890625, 4743.51318359375, 
    4693.23486328125, 4541.75048828125, 4595.9609375, 4739.77392578125, 
    4739.77392578125, 4941.40185546875, 4850.2900390625, 4973.033203125, 
    4884.119140625, 4680.42626953125, 4739.4521484375, 4588.32373046875, 
    4741.61865234375, 4276.41748046875, 1765.66845703125, -0, -0, -0, -0, 
    888.764831542969, 1440.57055664062, 1420.41052246094, 1308.09875488281, 
    1401.07348632812, 1759.77270507812, 2524.69189453125, 2724.66137695312, 
    2559.86596679688, 2596.80322265625, 3552.53198242188, 3694.46069335938, 
    3514.53442382812, 3982.24487304688, 4326.27490234375, 4821.6083984375, 
    4779.07571895829, 5021.10888671875, 5190.2021484375, 5279.1142578125, 
    5267.3056640625, 5380.2060546875, 5447.91064453125, 5414.7158203125, 
    5452.94970703125, 5288.201171875, 5247.45166015625, 4978.1376953125, 
    4977.318359375, 4715.31640625, 4715.31640625, 4255, 4345.37109375, 
    4345.37109375, 4690.06884765625, 5050.8427734375, 5050.8427734375, 
    5046.09716796875, 5083.7783203125, 5132.41162109375, 4992.9580078125, 
    5045.52880859375, 5045.52880859375, 5008.66259765625, 5198.9326171875, 
    5301.21923828125, 5264.1083984375, 5165.62451171875, 5167.36865234375, 
    5031.37451171875, 5226.81689453125, 5347.77783203125, 5330.63671875, 
    5016.52490234375, 5038.005859375, 4980.51416015625, 4908.0869140625, 
    4800.0302734375, 4817.49951171875, 4741.59912109375, 4696.0283203125, 
    4603.65185546875, 4502.8251953125, 4421.185546875, 4235.3974609375, 
    4033.23681640625, 4033.23681640625, 3987.8662109375, 3939.87866210938, 
    3666.841796875, 3233.7724609375, 3339.47192382812, 3350.44946289062, 
    3262.16259765625, 3066.64331054688, 2695.33227539062, 2662.02612304688, 
    2972.39501953125, 3095.21997070312, 3192.92431640625, 3334.51733398438, 
    3323.08154296875, 3526.533203125, 3506.61669921875, 3721.27612304688, 
    3729.39916992188, 3823.66577148438, 3869.82080078125, 4170, 4170, 
    4297.306640625, 4206.1083984375, 4209.60791015625, 4175, 4175, 4175, 
    4228.5361328125, 4108.044921875, 4175, 4025.4287109375, 3705.10009765625, 
    3907.53588867188, 4085.73364257812, 4335.14208984375, 4053.87622070312, 
    3426.97705078125, 3452.13110351562, 3286.33715820312, 3252.31713867188, 
    3162.25415039062, 2644.24951171875, 2724.3701171875, 2724.3701171875, 
    683.282409667969, -0, -0, -0, -0, -0, -0, -0, -0, 90, 90, 90, 90, 80, 
    110, 120, 1122.97009277344, 2498.4326171875, 3871.24682617188, 
    5339.12158203125, 5468.94482421875, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5355.458984375, 5278.95849609375, 5178.59423828125, 5158.427734375, 
    5203.0400390625, 5307.08544921875, 5348.134765625, 5285.8193359375, 
    5223.5244140625, 5318.3564453125, 5385.8193359375, 5473.69091796875, 
    5500, 5500, 5326.22412109375, 5300.810546875, 5184.2021484375, 
    4947.81787109375, 4888.2216796875, 4674.359375, 4602.4677734375, 
    4638.09033203125, 4501.17529296875, 4352.79052734375, 4179.638671875, 
    3997.66723632812, 3994.56909179688, 3989.6708984375, 3768.59912109375, 
    3699.28247070312, 3387.2978515625, 3314.40454101562, 2794.44604492188, 
    2551.75659179688, 3017.04833984375, 3261.50463867188, 3068.17724609375, 
    3096.03857421875, 3429.65991210938, 3561.74853515625, 3617.67358398438, 
    3616.92358398438, 3681.10888671875, 3681.10888671875, 3683.71557617188, 
    3722.0029296875, 3965.26538085938, 3889.18017578125, 3575.5576171875, 
    4278.58544921875, 4548.150390625, 4427.4912109375, 3902.515625, 
    3902.515625, 3855.0078125, 4225.23046875, 4387.0732421875, 
    4508.931640625, 4741.80615234375, 4746.6513671875, 4653.7080078125, 
    4699.7216796875, 4699.7216796875, 4663.91748046875, 4656.99072265625, 
    4505.78857421875, 4533.78564453125, 4315.1044921875, 4483.2998046875, 
    4725.3486328125, 4885.2861328125, 5027.7939453125, 5089.96435546875, 
    5500, 5500, 5500, 5500, 5275.9541015625, 5270.296875, 4739.34619140625, 
    4045.85375976562, 3749.66625976562, 2495.6123046875, 2102.31860351562, 
    2366.74951171875, 2376.2080078125, 1903.154296875, 1903.154296875, 
    1830.53381347656, 1349.80310058594, 1517.73693847656, 1652.23681640625, 
    1652.23681640625, 1504.39001464844, 1507.44494628906, 2158.93725585938, 
    2158.93725585938, 1303.64562988281, 995.814575195312, 2274.869140625, 
    3065.78548661781, 3365.74584960938, 3532.3720703125, 4046.8798828125, 
    4262.93017578125, 4419.18185522252, 4511.8134765625, 4630.58203125, 
    4703.26220703125, 4703.93896484375, 4532.01416015625, 4656.03662109375, 
    4640.16064453125, 4248.00927734375, 3598.24243164062, 2680.8271484375, 
    3206.044921875, 3387.2978515625, 3685.79858398438, 3451.85595703125, 
    3609.23754882812, 3672.345703125, 3577.20141601562, 3541.64819335938, 
    3546.8037109375, 3533.37231445312, 3416.09521484375, 3461.81225585938,
  3399.08178710938, 3454.22143554688, 3424.04614257812, 3408.71313476562, 
    3410.11669921875, 3397.8857421875, 3426.8076171875, 3413.08129882812, 
    3234.44067382812, 3204.49169921875, 3127.96630859375, 3047.92260742188, 
    3047.92260742188, 2923.28002929688, 2910.35009765625, 3043.72875976562, 
    3066.55712890625, 3259.44287109375, 3346.48852539062, 3637.16845703125, 
    3669.06127929688, 3629.14697265625, 3658.85522460938, 3630.224609375, 
    3646.02758789062, 3757.56494140625, 3945.54052734375, 4015.74584960938, 
    3991.27807617188, 4032.64477539062, 4032.64477539062, 4108.68896484375, 
    4172.1279296875, 4182.046875, 4253.7431640625, 4250.8486328125, 
    4187.087890625, 4320.99365234375, 4348.435546875, 4364.15185546875, 
    4439.78564453125, 4542.4658203125, 4520.63330078125, 4497.26953125, 
    4400.96484375, 4528.80322265625, 4628.779296875, 4691.8212890625, 
    4801.7734375, 4971.6181640625, 4712.27734375, 4648.6943359375, 
    4665.6328125, 4591.43017578125, 4605.33740234375, 4575.67578125, 
    4539.42333984375, 4533.9072265625, 4423.5146484375, 4643.71337890625, 
    4732.466796875, 4696.47021484375, 4632.1552734375, 4632.1552734375, 
    3925.75561523438, 2666, 2666, 2666, 3535, 4035, 4035, 4027.89575195312, 
    4652.0693359375, 4618.572265625, 4660.740234375, 4739.77392578125, 
    4739.77392578125, 4607.61572265625, 4850.2900390625, 4962.3154296875, 
    5015.52978515625, 4891.828125, 4765.8671875, 4765.77294921875, 
    4760.69677734375, 4276.41748046875, 3703.88037109375, 2003.99548339844, 
    -0, -0, -0, 130, 180, 659.17626953125, 737.6005859375, 741.584533691406, 
    971.206420898438, 1283.15771484375, 1354.75463867188, 1465.75073242188, 
    1102.48132324219, 901.071411132812, 814.165405273438, 413.3017578125, 
    874.808410644531, 2221.57763671875, 3387.2978515625, 4209.5869140625, 
    4548.44921875, 4896.85400390625, 5198.24462890625, 5156.83984375, 
    5252.78369140625, 5320.65869140625, 5373.5771484375, 5296.6337890625, 
    5128.52197265625, 5076.017578125, 4978.1376953125, 4668.08056640625, 
    4665, 5016.791015625, 4848.27001953125, 4792.25, 4257.06298828125, 
    4891.25830078125, 5059.1328125, 5059.1328125, 5054.42822265625, 
    5048.751953125, 5187.73583984375, 5197.46728515625, 5180.20361328125, 
    5103.91650390625, 5097.95703125, 5196.1328125, 5294.595703125, 
    5416.54443359375, 5385.98193359375, 5267.796875, 5161.73583984375, 
    5170.2587890625, 5345.08251953125, 5167.2490234375, 5016.52490234375, 
    5017.93798828125, 4935.02587890625, 4900.3232421875, 4975.76318359375, 
    5017.9638671875, 4896.86083984375, 4693.7724609375, 4688.3408203125, 
    4658.4873046875, 4490.412109375, 4395.72509765625, 4314.01416015625, 
    4242.62158203125, 3971.00048828125, 3988.46655273438, 3561.12744140625, 
    3538.32836914062, 3653.08081054688, 3528.13134765625, 3402.54565429688, 
    3198.19384765625, 2955.08422851562, 2788.45361328125, 2901.52954101562, 
    3082.51220703125, 3239.51611328125, 3104.583984375, 3274.64135742188, 
    3433.13061523438, 3591.99365234375, 3694.69970703125, 3790.57666015625, 
    3844.54614257812, 3857.3125, 4170, 4170, 4065.89147763595, 
    4205.1748046875, 4033.19677734375, 4194.27880859375, 4133.15185546875, 
    4311.0732421875, 4275.35986328125, 4264.5302734375, 4197.27880859375, 
    4034.73999023438, 3897.55419921875, 3775.71533203125, 3728.04833984375, 
    3663.77294921875, 3505.25732421875, 3400.14038085938, 2829.68188476562, 
    3134.134765625, 3277.83715820312, 3367.35034179688, 3355.1416015625, 
    2984.19580078125, 2984.19580078125, 1236.67016601562, 0, 0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 90, 90, 80, 110, 120, 1122.97009277344, 
    2136.69848632812, 3879.888671875, 5157.439453125, 5415.54931640625, 5500, 
    5500, 5500, 5500, 5500, 5380.69970703125, 5255.45263671875, 
    5192.724609375, 5056.724609375, 5064.88134765625, 5061.9375, 
    5104.21337890625, 5104.21337890625, 5110.0556640625, 5085.5556640625, 
    5089.466796875, 5234.1494140625, 5349.52490234375, 5337.36767578125, 
    5339.8251953125, 5313.57177734375, 5327.30810546875, 5245.6044921875, 
    5078.41162109375, 4947.81787109375, 4648.91162109375, 4582.46435546875, 
    4610.23095703125, 4427.603515625, 4474.0869140625, 4648.5546875, 
    4376.787109375, 4206.41015625, 3858.25756835938, 3814.27563476562, 
    3695.9169921875, 3545.07470703125, 3403.9658203125, 2965.18359375, 
    2966.25439453125, 3291.08862304688, 3596.46630859375, 3402.74243164062, 
    3476.4033203125, 3603.04736328125, 3639.8935546875, 3690.57177734375, 
    3676.1806640625, 3775.56762695312, 3721.27612304688, 3677.35571289062, 
    3317.25244140625, 3710.30322265625, 3889.18017578125, 3967.2138671875, 
    4048.25708007812, 4380.70654296875, 4394.4765625, 3834.08837890625, 
    3289.96850585938, 3855.0078125, 3855.0078125, 4361.83935546875, 
    4387.0732421875, 4666.8291015625, 4666.421875, 4666.421875, 
    4795.01904296875, 4840.6787109375, 4781.19287109375, 5064.81103515625, 
    4816.87109375, 4806.560546875, 4542.9052734375, 4559.63134765625, 
    4340.96728515625, 4763.1181640625, 4922.77734375, 4997.67822265625, 
    5089.96435546875, 5203.24658203125, 5500, 5500, 5500, 5473.08203125, 
    5152.6162109375, 4963.58251953125, 4728.04248046875, 4331.373046875, 
    3851.26879882812, 3626.03930664062, 2024.54443359375, 2070.14599609375, 
    1903.154296875, 2144.58056640625, 2246.56762695312, 2246.56762695312, 
    2223.48583984375, 2297.24096679688, 1612.21337890625, 1722.00354003906, 
    2060.16748046875, 2424.2744140625, 2354.11157226562, 2227.099609375, 
    2973.91674804688, 3257.98315429688, 3483.71728515625, 3566.9580078125, 
    3796.7060546875, 4246.0126953125, 4376.4208984375, 4530.83935546875, 
    4666.89599609375, 4696.82177734375, 4810.19384765625, 4854.6630859375, 
    4854.71142578125, 4850.05224609375, 4779.07571895829, 4524.33837890625, 
    4447.72314453125, 4074.40869140625, 3839.044921875, 3970.9638671875, 
    3904.83862304688, 3695.14477539062, 3647.60034179688, 3686.52416992188, 
    3450, 3547.18774414062, 3697.423828125, 3430.76684570312, 
    3423.64282226562, 3415.26489257812,
  3291.21728515625, 3157.23461914062, 3255.5478515625, 3218.28442382812, 
    3209.958984375, 3194.05590820312, 3173.02026367188, 3075.98071289062, 
    3047.27099609375, 2965.701171875, 2963.49169921875, 2819.91235351562, 
    2741.81176757812, 2910.29345703125, 3055.45263671875, 3173.53833007812, 
    3317.78564453125, 3387.2978515625, 3569.48876953125, 3655.71215820312, 
    3784.18530273438, 3774.3662109375, 3863.15356445312, 3790.15625, 
    3822.73901367188, 3930.33837890625, 3950.69799804688, 4068.73510742188, 
    4132.490234375, 4098.078125, 4141.20654296875, 4318.3994140625, 
    4311.705078125, 4327.25244140625, 4393.349609375, 4292.01611328125, 
    4253.4814453125, 4419.18185522252, 4498.576171875, 4495.1982421875, 
    4526.47119140625, 4587.16796875, 4573.31982421875, 4612.83935546875, 
    4603.70068359375, 4566.630859375, 4618.46923828125, 4779.07571895829, 
    4779.07571895829, 4841.79736328125, 4864.0244140625, 4909.92041015625, 
    4878.9228515625, 4836.54541015625, 4803.05908203125, 4688.2294921875, 
    4730.05908203125, 4722.5537109375, 4613.17626953125, 4577.55859375, 
    4577.55859375, 4709.38525390625, 4739.619140625, 4702.67529296875, 
    3539.6123046875, 1152.67797851562, -0, 80, 3041.84375, 3041.84375, 
    2879.25903320312, 4181.49072265625, 4671.01513671875, 4618.572265625, 
    4623.6884765625, 4694.58349609375, 4694.58349609375, 4566.21923828125, 
    4634.07177734375, 4962.3154296875, 5025.49560546875, 4966.6279296875, 
    4765.8671875, 4765.77294921875, 4004.74853515625, 4004.74853515625, 
    3703.88037109375, 2441.4501953125, 1134.22229003906, 140, -0, -0, -0, 
    150, 210, 210, 270.610395222517, 270.610395222517, 392.007965087891, 
    430.492309570312, 437.623107910156, 402.218902587891, 270.610395222517, 
    253.361404418945, 760.75927734375, 1136.10766601562, 1715.13916015625, 
    2073.80419921875, 2370.75122070312, 4000.76171875, 4108.53125, 
    4351.3623046875, 5090.65771484375, 5368.82421875, 5257.77490234375, 
    5185.01708984375, 5085.23583984375, 5108.86083984375, 4010, 
    4966.93017578125, 5124.36572265625, 4848.27001953125, 4956.529296875, 
    4972.77001953125, 4959.48388671875, 4989.10986328125, 5059.1328125, 
    5143.41858983545, 5205.52294921875, 5212.44921875, 5216.3046875, 
    5331.349609375, 5323.673828125, 5459.47802734375, 5242.6015625, 
    5205.0263671875, 5335.6904296875, 5409.42236328125, 5425.7802734375, 
    5435.62744140625, 5248.7744140625, 5454.52587890625, 5237.88720703125, 
    5247.04833984375, 4961.0478515625, 5083.66845703125, 5039.4140625, 
    5078.24462890625, 5037.45703125, 4997.23095703125, 4962.1484375, 
    4718.60107421875, 4728.3720703125, 4685.099609375, 4558.55712890625, 
    4395.44189453125, 4302.3681640625, 4132.82470703125, 3779.30615234375, 
    3668.66552734375, 3722.0439453125, 3924.7705078125, 3923.88232421875, 
    3670.671875, 3529.078125, 3274.93481445312, 3135.56176757812, 
    2877.77392578125, 2758.41088867188, 3077.21533203125, 3250.97729492188, 
    3192.70629882812, 3300.23364257812, 3475.99340820312, 3548.716796875, 
    3732.13549804688, 3794.9404296875, 3860.35205078125, 3987.15063476562, 
    4171.94677734375, 4251.8642578125, 4113.80908203125, 4190, 
    4234.27880859375, 4111.65869140625, 4181.595703125, 4289.54736328125, 
    4327.37890625, 4142.5, 4210.58154296875, 4034.73999023438, 
    3867.41259765625, 3534.04296875, 3503.7861328125, 3510.04711914062, 
    3289.05834960938, 3269.33422851562, 2832.4892578125, 3175.01220703125, 
    3363.57958984375, 3511.10009765625, 3572.921875, 3342.49438476562, 
    3342.49438476562, 2634.23681640625, 485, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 60, 60, 80, 90, 90, 522.4765625, 2010.9462890625, 3322.81298828125, 
    4726.79150390625, 5162.0576171875, 5500, 5500, 5500, 5500, 
    5399.44677734375, 5372.7802734375, 5336.1474609375, 5214.15966796875, 
    5197.818359375, 5095.9970703125, 5173.06103515625, 5186.2626953125, 
    5171.693359375, 5177.837890625, 5190.32763671875, 5175.8603515625, 
    5241.77587890625, 5307.80712890625, 5210.4208984375, 5143.41858983545, 
    5078.19580078125, 5022.384765625, 4891.39599609375, 4917.494140625, 
    4696.36669921875, 4561.595703125, 4581.75439453125, 4603.2080078125, 
    4614.98681640625, 4619.6103515625, 4532.4775390625, 4376.787109375, 
    4082.91162109375, 3797.65307617188, 3721.70751953125, 3650.97338867188, 
    3405.32958984375, 3147.9970703125, 2572.68408203125, 2966.25439453125, 
    3291.08862304688, 3388.35888671875, 3653.84741210938, 3606.32397460938, 
    3624.26879882812, 3709.21142578125, 3693.26733398438, 3837.31005859375, 
    4128.744140625, 4235.78466796875, 3361.76538085938, 3593.50366210938, 
    3593.50366210938, 2382.77612304688, 3967.2138671875, 4028.61840820312, 
    4240.82666015625, 4240.82666015625, 4364.29052734375, 4602.55517578125, 
    4555.08837890625, 4077.81030273438, 3253.61059570312, 4181.05224609375, 
    4119.00341796875, 4421.01416015625, 4695.58447265625, 4783.1904296875, 
    4899.3564453125, 4971.8212890625, 5009.2060546875, 4864.72900390625, 
    4837.1826171875, 4789.724609375, 4864.67822265625, 4992.88525390625, 
    4880.53466796875, 4779.07571895829, 4849.5947265625, 5131.31640625, 
    5055.005859375, 5224.67529296875, 5217.69091796875, 5436.61083984375, 
    5407.7646484375, 5425.66455078125, 5294.4111328125, 4728.04248046875, 
    4728.04248046875, 4075.23559570312, 4123.96875, 3250.88500976562, 
    3163.31860351562, 2638.57250976562, 2577.83276367188, 2525.603515625, 
    2314.4853515625, 2994.09301757812, 2805.74755859375, 2615.8310546875, 
    2615.8310546875, 2605.3603515625, 2427.81079101562, 2354.11157226562, 
    2227.099609375, 2798.43237304688, 3221.77001953125, 3496.48022460938, 
    3809.60205078125, 4089.03515625, 4308.9853515625, 4578.0224609375, 
    4686.986328125, 4646.4375, 4881.41796875, 4988.44287109375, 
    5101.41845703125, 5055.72802734375, 4802.48388671875, 4799.09716796875, 
    4664.95263671875, 4475.1337890625, 4306.02587890625, 4138.74609375, 
    3965.6318359375, 4008.15551757812, 3869.56787109375, 3734.9228515625, 
    3721.27612304688, 3453.37768554688, 3302.36352539062, 3142.32861328125, 
    3286.23754882812, 3297.39990234375, 3291.06787109375,
  2942.03344726562, 2775.91137695312, 2739.34545898438, 2801.55517578125, 
    2992.40454101562, 2992.40454101562, 2858.6611328125, 2855.83642578125, 
    2758.41088867188, 2724.93725585938, 2731.2470703125, 2921.61596679688, 
    3154.46142578125, 3178.037109375, 3218.84838867188, 3353.9501953125, 
    3406.48657226562, 3546.63549804688, 3632.86645507812, 3695.17163085938, 
    3848.74951171875, 3992.95092773438, 3866.11865234375, 3886.87353515625, 
    3947.9111328125, 3921.76733398438, 4116.8720703125, 4156.8193359375, 
    4300.8232421875, 4172.06494140625, 4314.6318359375, 4324.77978515625, 
    4324.86328125, 4366.92822265625, 4357.7294921875, 4451.1416015625, 
    4437.7578125, 4574.62548828125, 4595.94775390625, 4577.154296875, 
    4687.20458984375, 4644.53759765625, 4619.18701171875, 4639.40234375, 
    4728.30224609375, 4728.30224609375, 4779.72021484375, 4956.75537109375, 
    4906.037109375, 5047.61572265625, 4968.3125, 5040.3525390625, 
    5071.5283203125, 4972.55615234375, 4903.28466796875, 4908.79638671875, 
    4862.5859375, 4870.38232421875, 4674.13916015625, 4675, 4681.41650390625, 
    4681.41650390625, 4681.41650390625, 4465.36083984375, 2155.33349609375, 
    -0, -0, -0, 882.829711914062, 3643.8193359375, 4298.00732421875, 
    4454.9990234375, 4664.837890625, 4681.298828125, 4552.71044921875, 
    4568.4990234375, 4698.9228515625, 4566.21923828125, 4613.35546875, 
    4784.53076171875, 4987.8974609375, 4959.57568359375, 4881.6787109375, 
    4626.802734375, 4128.40380859375, 4402.9521484375, 3697.78662109375, 
    2191.85384798669, 1134.22229003906, 942.839303029559, 370.154968261719, 
    -0, -0, -0, 210, 210, 1777.81384277344, 2014.4833984375, 
    2016.99096679688, 1872.99035644531, 1896.08569335938, 1777.65539550781, 
    1823.9228515625, 2411.30908203125, 2338.46020507812, 2237.86401367188, 
    1985.20458984375, 1788.74865722656, 1906.54235839844, 2434.6416015625, 
    2986.03173828125, 2775.705078125, 4679.21142578125, 4894.58154296875, 
    4910.8779296875, 5067.11083984375, 5056.34423828125, 4216.89208984375, 
    5084.23486328125, 5084.23486328125, 5006.31396484375, 4904.0283203125, 
    4828.8515625, 4819.2021484375, 5011.34326171875, 4989.10986328125, 
    5117.8037109375, 5201.02001953125, 5244.93408203125, 5148.84912109375, 
    5206.62841796875, 5350.43896484375, 5316.87646484375, 5500, 5500, 
    5476.4169921875, 5485.9013671875, 5393.58837890625, 5309.6181640625, 
    5500, 5500, 5273.9599609375, 5222.87548828125, 5193.8583984375, 
    5063.75439453125, 4999.72314453125, 5048.50537109375, 5039.4140625, 
    5010.09912109375, 5025.890625, 4833.93408203125, 4708.93115234375, 
    4620.1220703125, 4603.2802734375, 4532.13671875, 4436.13427734375, 
    4306.9072265625, 4117.86083984375, 3935.38159179688, 4033.26635742188, 
    4018.64526367188, 3954.41528320312, 3829.54321289062, 3670.671875, 
    3530.80786132812, 3274.93481445312, 3162.31127929688, 2825.37158203125, 
    2589.93969726562, 2928.61328125, 3198.4091796875, 3186.44116210938, 
    3272.9560546875, 3375.87524414062, 3524.68920898438, 3757.7197265625, 
    3897.712890625, 3918.00366210938, 4031.18774414062, 4171.94677734375, 
    4187.08349609375, 4260.33837890625, 4190, 4228.87939453125, 4336.4765625, 
    4277.08740234375, 4180.068359375, 4155.79443359375, 3973.05981445312, 
    3813.73022460938, 3800.49658203125, 3924.95190429688, 3680.59912109375, 
    3480.787109375, 3357.61694335938, 3017.44262695312, 2741.85302734375, 
    2956.18115234375, 3369.53466796875, 3363.57958984375, 3407.52612304688, 
    3535.3828125, 3342.49438476562, 3361.71337890625, 3361.71337890625, 485, 
    0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 80, 80, 90, 90, 
    596.518188476562, 1808.90026855469, 3654.84838867188, 4812.62890625, 
    5359.443359375, 5500, 5500, 5500, 5500, 5500, 5500, 5275.3125, 
    5214.2177734375, 5095.9970703125, 5143.41858983545, 5192.21533203125, 
    5185.12841796875, 5157.16357421875, 5166.34033203125, 5173.63623046875, 
    5175.03076171875, 5198.900390625, 5198.125, 5114.455078125, 5006.9453125, 
    5006.9453125, 4954.8818359375, 4621.41259765625, 4438.84912109375, 
    4518.8564453125, 4465.99560546875, 4513.2158203125, 4580.9296875, 
    4489.99267578125, 4383.6416015625, 4255.38525390625, 3901.92016601562, 
    3724.61474609375, 3524.23461914062, 3485.3125, 3234.58959960938, 
    3088.15405273438, 2446.94750976562, 2802.7392578125, 3144.19506835938, 
    3142.52075195312, 3322.37329101562, 3606.32397460938, 3697.61840820312, 
    3594.7216796875, 3697.20825195312, 3793.57299804688, 4115.92431640625, 
    4258.03857421875, 4101.1005859375, 4218.10595703125, 4268.4970703125, 
    1636.6259765625, 1737.7939453125, 2784.06396484375, 3304.1884765625, 
    3670.66259765625, 4354.42529296875, 4705.2236328125, 4748.82177734375, 
    4748.82177734375, 4748.82177734375, 4548.154296875, 4219.72216796875, 
    3614.55932617188, 3907.75610351562, 4577.08056640625, 4671.72412109375, 
    5081.4326171875, 4948.98828125, 4931.6123046875, 4931.6123046875, 
    4831.7685546875, 5019.83935546875, 5112.07470703125, 5096.87255859375, 
    4556.38525390625, 3785.95532226562, 3850.24169921875, 4291.73828125, 
    4555.56298828125, 4672.20556640625, 4693.7841796875, 5041.40625, 
    5239.21142578125, 5198.5009765625, 4880.2734375, 4811.57275390625, 
    4614.48681640625, 4122.31201171875, 4122.31201171875, 3816.13330078125, 
    3100.46020507812, 2837.47973632812, 2606.71313476562, 2314.4853515625, 
    2932.90966796875, 2805.74755859375, 3134.95385742188, 3339.62939453125, 
    3105.31201171875, 2996.814453125, 2958.73999023438, 2851.35888671875, 
    3081.66040039062, 3651.76489257812, 3496.48022460938, 3918.96118164062, 
    4199.39453125, 4401.6708984375, 4466.99755859375, 4668.505859375, 
    4849.76123046875, 4835.953125, 4941.52294921875, 5026.298828125, 
    5026.298828125, 4992.5546875, 4943.96240234375, 4704.34521484375, 
    4332.77197265625, 4346.02685546875, 4199.31884765625, 4164.94970703125, 
    4083.89916992188, 3943.11743164062, 3983.01196289062, 3840.1025390625, 
    3647.81811523438, 3309.96166992188, 3132.54028320312, 3065.78548661781, 
    3044.26000976562, 2976.55688476562,
  2970.96215820312, 2658.537109375, 2768.73168945312, 3065.78548661781, 
    3174.611328125, 3217.99096679688, 2688.533203125, 2679.87426757812, 
    2651.22485351562, 2626.11352539062, 2933.23413085938, 3127.88330078125, 
    3201.748046875, 3341.95483398438, 3399.33374023438, 3533.45556640625, 
    3535.67944335938, 3664.74340820312, 3808.662109375, 3996.94921875, 
    3975.85375976562, 4116.7626953125, 4246.375, 4135.451171875, 
    4031.81469726562, 4123.09375, 4301.2333984375, 4187.48486328125, 
    4384.666015625, 4398.25390625, 4377.2685546875, 4395.8935546875, 
    4449.94873046875, 4454.1669921875, 4475.77099609375, 4523.841796875, 
    4514.6650390625, 4552.1650390625, 4653.466796875, 4653.466796875, 
    4851.17822265625, 4858.060546875, 4701.59814453125, 4990.34912109375, 
    4945.40283203125, 4916.47265625, 4926.02734375, 5008.6201171875, 
    5069.12890625, 5189.91064453125, 5357.81640625, 5179.90673828125, 
    5077.4599609375, 5118.65576171875, 5044.0751953125, 4996.62353515625, 
    4988.5859375, 4988.3564453125, 4674.13916015625, 4961.4375, 
    5098.5244140625, 4681.41650390625, 4538.91943359375, 3256.49829101562, 
    370.154968261719, -0, -0, -0, 270.610395222517, 3933.146484375, 
    4621.54736328125, 4749.19189453125, 4615.11279296875, 4738.75830078125, 
    4744.4013671875, 4419.18185522252, 4441.45458984375, 4530.33544921875, 
    4584.935546875, 4779.07571895829, 4900.00537109375, 4809.1005859375, 
    4840.72705078125, 4688.6962890625, 4128.40380859375, 4240.78369140625, 
    3479.49560546875, 1434.54553222656, 1034.98815917969, 948.688354492188, 
    547.00830078125, 180, -0, -0, 140, 190, 1844.57434082031, 
    2014.4833984375, 2856.39697265625, 2773.634765625, 2645.326171875, 
    2601.70458984375, 3038.89672851562, 3038.89672851562, 3101.87426757812, 
    3221.37255859375, 3196.3154296875, 3640.3505859375, 3663.09399414062, 
    3908.72705078125, 4316.28564453125, 4129.01953125, 4676.6162109375, 
    4885.736328125, 5053.16943359375, 3657.29223632812, 4923.61572265625, 
    5009.494140625, 5182.806640625, 5229.443359375, 5006.31396484375, 
    5027.48193359375, 4942.626953125, 4887.35693359375, 4933.6748046875, 
    4964.92138671875, 5052.91748046875, 5099.552734375, 5148.44287109375, 
    5143.41858983545, 5254.47509765625, 5363.650390625, 5479.42919921875, 
    5500, 5500, 5500, 5475.62451171875, 5349.7734375, 5500, 5392.9814453125, 
    5280.6005859375, 5195.1796875, 5098.84326171875, 5098.84326171875, 
    5079.69921875, 5001.3408203125, 5075.49609375, 5121.0830078125, 
    4997.19580078125, 4946.4033203125, 4862.95166015625, 4718.18310546875, 
    4674.5634765625, 4576.076171875, 4546.9052734375, 4437.173828125, 
    4122.2451171875, 4163.63818359375, 4115.26806640625, 4079.25219726562, 
    4091.525390625, 3869.08032226562, 3777.81420898438, 3611.10717773438, 
    3420.78491210938, 3132.64184570312, 2974.66235351562, 2864.3359375, 
    2708.31225585938, 2881.23046875, 3140.85986328125, 3314.27880859375, 
    3476.74780273438, 3538.52221679688, 3671.59619140625, 3595.49926757812, 
    3863.34497070312, 3991.7412109375, 4031.18774414062, 4065.89147763595, 
    4187.08349609375, 4187.08349609375, 3999.43823242188, 3868.17822265625, 
    3740.50341796875, 3818.10131835938, 3667.58276367188, 3538.36059570312, 
    3442.17016601562, 3349.72875976562, 3171.37036132812, 3680.59912109375, 
    3680.59912109375, 3572.67919921875, 3572.67919921875, 3292.01684570312, 
    3418.77685546875, 3596.82397460938, 3652.15356445312, 3548.5322265625, 
    3612.67211914062, 3675.40747070312, 3675.40747070312, 3674.11352539062, 
    3674.11352539062, 542.932983398438, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    40, 40, 40, 60, 70, 80, 90, 339.273620605469, 1745.70373535156, 
    4300.97119140625, 4830.23095703125, 5400.59765625, 5495.1015625, 5500, 
    5500, 5500, 5500, 5341.103515625, 5124.8720703125, 5115.12744140625, 
    5117.18798828125, 5168.02099609375, 5185.0927734375, 5179.86669921875, 
    5197.50244140625, 5208.912109375, 5211.2734375, 5230.36572265625, 
    5227.11865234375, 5038.89697265625, 4961.64599609375, 4903.73291015625, 
    4872.14208984375, 4715.8037109375, 4695.669921875, 4654.21142578125, 
    4487.1728515625, 4476.92431640625, 4470.94775390625, 4354.8525390625, 
    4219.82421875, 4023.24462890625, 3905.21557617188, 3668.45703125, 
    3570.74438476562, 3472.53662109375, 3331.32739257812, 2759.57275390625, 
    2644.42260742188, 2945.39038085938, 3129.572265625, 3088.63623046875, 
    3297.56811523438, 3569.83813476562, 3594.7216796875, 3594.7216796875, 
    3697.20825195312, 3762.69116210938, 3951.19506835938, 4121.62109375, 
    4340.69287109375, 4219.65869140625, 4095.0546875, 3680.30981445312, 
    3121.54052734375, 3247.27685546875, 3827.39721679688, 4050.88403320312, 
    4530.392578125, 4742.755859375, 4802.2919921875, 4779.07571895829, 
    4878.43603515625, 4735.599609375, 4660.96728515625, 4621.05419921875, 
    4764.3017578125, 3602.04345703125, 4125.82861328125, 4514.09375, 
    4930.89111328125, 4931.6123046875, 4962.6435546875, 4831.7685546875, 
    5087.85107421875, 5069.62646484375, 5104.171875, 4970.2578125, 
    4200.85546875, 3215.59692382812, 2772.11254882812, 3080.88159179688, 
    3085.01025390625, 4139.6640625, 4914.85986328125, 4974.69775390625, 
    4921.220703125, 4880.2734375, 4857.06103515625, 4902.814453125, 
    4684.9404296875, 4228.005859375, 3864.998046875, 3559.89892578125, 
    3270.00732421875, 2808.74658203125, 2222.37451171875, 2358.84008789062, 
    2358.84008789062, 3374.48901367188, 3147.4931640625, 3130.73266601562, 
    2996.814453125, 3224.4140625, 3152.22509765625, 3425.57739257812, 
    3425.57739257812, 3387.2978515625, 4211.671875, 4347.70849609375, 
    4581.685546875, 4676.6748046875, 4797.35888671875, 4951.8818359375, 
    4926.1376953125, 4926.81396484375, 5029.41015625, 5123.44970703125, 
    5058.1064453125, 4873.130859375, 4619.57177734375, 4333.93359375, 
    4234.541015625, 4120.7177734375, 4086.064453125, 4065.89147763595, 
    4065.89147763595, 4079.25048828125, 3770.83471679688, 3619.06884765625, 
    3309.96166992188, 3203.58349609375, 3065.78548661781, 2901.37670898438, 
    2925,
  3115.56909179688, 3116.8642578125, 3094.83081054688, 3222.8017578125, 
    3299.34033203125, 3300.4150390625, 3102.8369140625, 2957.84375, 
    3025.51538085938, 3135.74877929688, 3198.10888671875, 3221.58544921875, 
    3342.50146484375, 3459.11669921875, 3533.880859375, 3652.73046875, 
    3771.462890625, 3868.81567382812, 3930.93627929688, 3930.93627929688, 
    3904.50268554688, 4275.7080078125, 4387.58447265625, 4328.45751953125, 
    4179.9345703125, 4356.3359375, 4360.92822265625, 4419.18185522252, 
    4446.17626953125, 4407.95556640625, 4545, 4545, 4572.6494140625, 
    4631.064453125, 4618.3671875, 4706.1357421875, 4699.87451171875, 
    4655.54443359375, 4851.54052734375, 4970.16162109375, 4792.31591796875, 
    4927.912109375, 4907.38232421875, 5171.673828125, 5154.04736328125, 
    5077.26806640625, 5098.38525390625, 5125.67724609375, 5231.796875, 
    5366.5712890625, 5311.97509765625, 5373.7685546875, 5379.48291015625, 
    5282.02392578125, 5264.23779296875, 5248.96044921875, 5205.15869140625, 
    5126.65576171875, 4880.68212890625, 4961.4375, 5019.4482421875, 
    4601.67822265625, 3400.27709960938, 479.242370605469, 60, 50, 50, 40, 80, 
    4025.00317382812, 4510.787109375, 4614.83984375, 4741.0908203125, 4690, 
    4644.13525390625, 4580, 4546.75341796875, 4591.1650390625, 4887.484375, 
    4923.31982421875, 4779.5908203125, 4728.42822265625, 4674.599609375, 
    4132.4130859375, 3664.41821289062, 3664.41821289062, 3027.25561523438, 
    1112.18237304688, 942.839303029559, 893.754638671875, 619.127075195312, 
    370.154968261719, 50, 50, -0, -0, -0, 1786.34680175781, 2773.634765625, 
    2938.23657226562, 2741.25561523438, 3308.3388671875, 3664.04272460938, 
    4078.0576171875, 4291.2783203125, 3888.29125976562, 4283.30615234375, 
    4396.34912109375, 4396.34912109375, 4319.9345703125, 4378.83837890625, 
    4378.83837890625, 4676.6162109375, 4676.6162109375, 3473.3837890625, 
    4881.76171875, 5064.37451171875, 5095.52392578125, 5320.49609375, 
    5154.068359375, 4993.72412109375, 4860.7734375, 4779.07571895829, 
    4814.72509765625, 4879.8076171875, 5016.2861328125, 4911.40966796875, 
    5017.5908203125, 5009.36962890625, 5186.53857421875, 5253.26708984375, 
    5464.5732421875, 5470.4775390625, 5500, 5431.43359375, 5400.11572265625, 
    5277.97119140625, 5500, 5410.10888671875, 5337.36962890625, 
    5425.86572265625, 5167.13623046875, 5037.0546875, 5058.02978515625, 
    5058.02978515625, 4973.93994140625, 4954.35205078125, 4993.1572265625, 
    5028.14794921875, 4903.873046875, 4801.86669921875, 4718.18310546875, 
    4568.79443359375, 4543.96630859375, 4386.21240234375, 4337.80908203125, 
    4087.73071289062, 4042.986328125, 4201.10888671875, 4258.240234375, 
    4314.2548828125, 4187.9716796875, 3915.51806640625, 3709.39306640625, 
    3507.54028320312, 3234.44018554688, 3104.09130859375, 3016.23901367188, 
    2583.14282226562, 2946.71752929688, 3103.29663085938, 3398.26953125, 
    3583.38110351562, 3721.27612304688, 3724.79321289062, 3777.2900390625, 
    3901.65380859375, 3971.65356445312, 3984.60302734375, 4174.50439453125, 
    4271.38916015625, 4315.8056640625, 3929.79614257812, 3747.1943359375, 
    3647.58813476562, 3623.6943359375, 3437.81860351562, 3169.37548828125, 
    2936.06567382812, 3204.09106445312, 3448.48364257812, 3518.89404296875, 
    3563.5283203125, 3684.62036132812, 3693.46508789062, 3683.15112304688, 
    3909.64819335938, 3787.59008789062, 4039.31616210938, 4219.07373046875, 
    4091.697265625, 3801.744140625, 3721.27612304688, 3957.07104492188, 
    3994.77978515625, 1243.64855957031, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 40, 60, 80, 90, 100, 520.021118164062, 1712.64733886719, 
    4181.93896484375, 5083.71337890625, 5393.54638671875, 5500, 
    5471.20458984375, 5489.9306640625, 5401.7197265625, 5253.080078125, 
    5169.513671875, 5117.5322265625, 5106.82958984375, 5131.17041015625, 
    5159.70556640625, 5176.3525390625, 5183.1064453125, 5192.33447265625, 
    5190.19189453125, 5270.35888671875, 5182.03857421875, 4978.64306640625, 
    5023.7685546875, 5018.8486328125, 4924.39501953125, 4715.8037109375, 
    4695.669921875, 4553.45458984375, 4339.98779296875, 4304.81591796875, 
    4327.3369140625, 4223.7978515625, 4128.01806640625, 3992.248046875, 
    3964.97534179688, 3853.66796875, 3535.99267578125, 3311.5, 
    3187.80786132812, 2966.14086914062, 2697.26782226562, 3016.26293945312, 
    3195.73486328125, 3141.228515625, 3217.02758789062, 3169.82348632812, 
    3223.51098632812, 3548.75048828125, 3447.69360351562, 3651.18188476562, 
    3420.54370117188, 3471.63061523438, 4100.5009765625, 4218.80517578125, 
    4374.93603515625, 4647.89208984375, 4675.3857421875, 4564.9560546875, 
    4723.57666015625, 4721.64990234375, 4819.21337890625, 5008.92431640625, 
    5090.69970703125, 5090.69970703125, 5064.41259765625, 4880.85693359375, 
    4789.69287109375, 4644.99267578125, 4710.55126953125, 4609.09521484375, 
    3728.9345703125, 1974.00964355469, 4097.47412109375, 4897.8681640625, 
    4948.1796875, 4948.6162109375, 4997.98583984375, 4987.35791015625, 
    5126.14794921875, 5126.14794921875, 4533.2783203125, 3492.87548828125, 
    2588.72387695312, 2453.1865234375, 2685.57836914062, 3602.20581054688, 
    4419.18185522252, 4518.44775390625, 4490.4423828125, 4284.39013671875, 
    4857.06103515625, 4934.78466796875, 4847.4150390625, 4585.26171875, 
    4214.9599609375, 4204.5107421875, 3799.9375, 3513.435546875, 
    2698.94946289062, 2171.16381835938, 2640.79760742188, 2640.79760742188, 
    2335.7890625, 2871.291015625, 2898.54150390625, 3109.55859375, 
    3315.10791015625, 3425.57739257812, 3782.4453125, 4046.8466796875, 
    4065.89147763595, 4303.0244140625, 4479.18701171875, 4752.51318359375, 
    4894.28466796875, 5060.38623046875, 5206.4228515625, 5202.4736328125, 
    5160.17529296875, 5133.11328125, 5072.8173828125, 4884.85107421875, 
    4524.708984375, 4313.23388671875, 4233.125, 4055.1533203125, 
    4055.1533203125, 4039.30322265625, 4171.20361328125, 4113.1455078125, 
    3871.60791015625, 3709.50512695312, 3603.9287109375, 3046.021484375, 
    2758.41088867188, 2784.79956054688, 3023.21948242188,
  3313.30004882812, 3345.40698242188, 3388.0244140625, 3422.93310546875, 
    3481.96655273438, 3509.23022460938, 3567.09545898438, 3576.98803710938, 
    3391.13159179688, 3424.44775390625, 3462.73657226562, 3358.01489257812, 
    3483.94604492188, 3553.01879882812, 3695.80688476562, 3760.37182617188, 
    3832.48315429688, 3926.15283203125, 4158.49462890625, 4233.4384765625, 
    4263.84912109375, 4226.9423828125, 4498.69140625, 4474.3486328125, 
    4482.05224609375, 4616.70458984375, 4524.19482421875, 4462.23388671875, 
    4419.18185522252, 4407.95556640625, 4596.82421875, 4598.37158203125, 
    4546.16357421875, 4680.5703125, 4732.13134765625, 4857.515625, 
    4824.73583984375, 4819.54638671875, 4845.31884765625, 4875.8193359375, 
    4904.36328125, 4820.16162109375, 5086.2275390625, 5322.69677734375, 
    5267.021484375, 5086.44677734375, 5130.19921875, 5242.0234375, 
    5263.88671875, 5367.4140625, 5464.8447265625, 5500, 5500, 5500, 5500, 
    5458.5595703125, 5353.2705078125, 5367.3662109375, 5012.404296875, 
    5122.134765625, 4353.25537109375, 3141.50341796875, 1611.14965820312, 90, 
    60, 50, 50, 40, 80, 3748.53369140625, 4472.69189453125, 4606.96142578125, 
    4704.06884765625, 4690, 4540, 4622.81103515625, 4580.52392578125, 
    4802.482421875, 4959.1396484375, 4903.8251953125, 4869.98974609375, 
    4664.31396484375, 4573.29833984375, 2576.59057617188, 2597.77368164062, 
    2553.662109375, 2553.662109375, 1062.74584960938, 638.99169921875, 
    619.127075195312, 775.971252441406, 683.282409667969, 200, 130, -0, -0, 
    -0, 180, 1841.78845214844, 3302.06396484375, 3344.36596679688, 
    3344.36596679688, 3864.1962890625, 4089.44506835938, 4678.48583984375, 
    4976.93115234375, 4852.45361328125, 4752.3896484375, 4612.80908203125, 
    4584.31982421875, 4635.76123046875, 4378.83837890625, 3959.21240234375, 
    3858.51538085938, 5094.5546875, 4881.76171875, 5064.37451171875, 
    5095.52392578125, 5095.52392578125, 5000.72900390625, 4726.904296875, 
    4755.29638671875, 4768.953125, 4768.953125, 4860.2705078125, 
    4857.88134765625, 4932.037109375, 5010.77099609375, 5143.41858983545, 
    5262.89306640625, 5431.83642578125, 5480.92431640625, 5463.5615234375, 
    5457.8154296875, 5382.24169921875, 5265.28857421875, 5500, 
    5316.28955078125, 5265.302734375, 5347.73095703125, 5168.21044921875, 
    4968.71826171875, 5037.0546875, 5041.46337890625, 5041.46337890625, 
    5028.72509765625, 4878.93359375, 5045.4736328125, 5007.08740234375, 
    4827.7802734375, 4609.76318359375, 4531.62109375, 4540.91357421875, 
    4531.45947265625, 4386.21240234375, 4351.009765625, 4198.8515625, 
    4224.98046875, 4311.13037109375, 4293.060546875, 4242.5205078125, 
    4154.5146484375, 3970.90747070312, 3709.39306640625, 3554.07421875, 
    3288.53662109375, 3190.31640625, 3008.55249023438, 2468.24829101562, 
    2897.65185546875, 3184.86206054688, 3393.6259765625, 3548.49975585938, 
    3721.27612304688, 3771.576171875, 3858.80493164062, 3875.92553710938, 
    3995.75610351562, 3984.60302734375, 4101.27880859375, 4271.38916015625, 
    4333.09033203125, 3709.1953125, 3644.75317382812, 3477.75146484375, 
    3318.5888671875, 3212.98803710938, 3211.23193359375, 3086.28100585938, 
    3204.09106445312, 3392.04736328125, 3583.20483398438, 3651.34521484375, 
    3684.62036132812, 4000.61743164062, 4000.61743164062, 3925.3466796875, 
    3787.59008789062, 3896.07275390625, 4065.89147763595, 4101.73779296875, 
    4103.48779296875, 3953.4609375, 3966.3740234375, 3966.3740234375, 
    1873.88439941406, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 
    60, 70, 90, 100, 761.006896972656, 2319.07202148438, 4493.56884765625, 
    4925.96533203125, 5295.6513671875, 5419.34228515625, 5376.62109375, 
    5371.3896484375, 5286.01025390625, 5193.791015625, 5168.92919921875, 
    5117.20556640625, 5102.19580078125, 5104.830078125, 5112.36962890625, 
    5123.24169921875, 5143.41858983545, 5183.99609375, 5167.2626953125, 
    5009.99755859375, 4938.85302734375, 5009.732421875, 4995.6748046875, 
    4836.7119140625, 4715.8037109375, 4689.9951171875, 4510.865234375, 
    4337.8193359375, 4246.98828125, 4234.1982421875, 4132.99267578125, 
    3968.52954101562, 4001.66870117188, 3993.64111328125, 3923.02001953125, 
    3745.65942382812, 3497.52563476562, 3211.97216796875, 2864.01513671875, 
    2591.39721679688, 2645.767578125, 2965.51147460938, 3106.59375, 
    3192.6591796875, 3169.82348632812, 3211.77075195312, 3070.12915039062, 
    3144.857421875, 3046.3916015625, 1242.09790039062, 3337.2939453125, 
    4183.50927734375, 4341.826171875, 4585.45166015625, 4745.26708984375, 
    4948.23681640625, 5090.63916015625, 5015.85009765625, 4999.08984375, 
    5071.44287109375, 5095.67822265625, 5111.65283203125, 5359.4345703125, 
    5332.271484375, 5171.3095703125, 4974.40380859375, 4779.07571895829, 
    4995.55908203125, 4720.880859375, 3728.9345703125, 4722.2587890625, 
    4827.1171875, 4913.44775390625, 4911.62109375, 5005.42041015625, 
    4791.31103515625, 5091.92724609375, 5126.14794921875, 5126.14794921875, 
    5009.75146484375, 3477.67919921875, 3555, 2673.10278320312, 
    3108.55200195312, 3934.65405273438, 4179.21142578125, 4179.21142578125, 
    3848.00390625, 4026.42358398438, 3977.04125976562, 4779.07571895829, 
    5409.80419921875, 5177.09326171875, 4848.76708984375, 4921.05029296875, 
    4391.00927734375, 3835.21240234375, 3123.01220703125, 2870.72314453125, 
    2640.79760742188, 2897.68676757812, 2938.20874023438, 2589.45874023438, 
    2439.86206054688, 3004.84228515625, 3315.10791015625, 3328.66381835938, 
    3782.4453125, 4046.8466796875, 4101.0322265625, 4152.27001953125, 
    4529.8857421875, 4752.51318359375, 5057.5966796875, 5203.130859375, 
    5323.3662109375, 5496.7099609375, 5313.29638671875, 5133.11328125, 
    4997.7890625, 4697.8603515625, 4648.66796875, 4383.7021484375, 
    4211.65771484375, 4155.19189453125, 4200.4326171875, 4186.37890625, 
    4287.54248046875, 4090.73583984375, 4079.1669921875, 3976.33325195312, 
    3603.9287109375, 3046.021484375, 1935.31774902344, 2355.59399414062, 
    3146.70703125,
  3341.484375, 3519.38818359375, 3514.76782226562, 3585.48583984375, 
    3587.42895507812, 3630.13427734375, 3650.62280273438, 3567.68994140625, 
    3591.0810546875, 3559.59521484375, 3635.607421875, 3635.607421875, 
    3631.51293945312, 3737.83081054688, 3744.59375, 3961.31420898438, 
    4065.89147763595, 4093.3134765625, 4275.5693359375, 4287.62548828125, 
    4384.43603515625, 4473.18798828125, 4603.37109375, 4546.85009765625, 
    4653.41650390625, 4653.41650390625, 4632.9013671875, 4656.74658203125, 
    4561.7138671875, 4565, 4565, 4568.43310546875, 4449.0009765625, 
    4352.20654296875, 4785.04443359375, 4827.82861328125, 5061.50634765625, 
    5039.064453125, 5025.57275390625, 4991.2490234375, 4957.943359375, 
    5014.7080078125, 5086.2275390625, 5285.62890625, 5359.70556640625, 
    5143.41858983545, 5114.21142578125, 5377.90478515625, 5488.07861328125, 
    5500, 5500, 5500, 5500, 5500, 5500, 5494.78955078125, 5500, 
    5498.07666015625, 5012.404296875, 3681.96020507812, 1596.55859375, 90, 
    40, -0, -0, 0, -0, 40, 80, 1770.14233398438, 4433.19384765625, 
    4555.6298828125, 4546.666015625, 4690.14013671875, 4540, 4541.4228515625, 
    4580.52392578125, 4907.5048828125, 4779.07571895829, 4732.25634765625, 
    4925.330078125, 4862.89013671875, 4761.31103515625, 2576.59057617188, 
    2313.22021484375, 2054.05590820312, 2157.36108398438, 742.064331054688, 
    524.6259765625, 534.035461425781, 753.9580078125, 1008.91186523438, 
    1008.91186523438, 282.838745117188, 150, -0, -0, -0, 294.462890625, 
    3302.06396484375, 3348.65063476562, 3348.65063476562, 3800.14184570312, 
    4287.95068359375, 4856.2421875, 5180.64990234375, 5245.7001953125, 
    5099.16943359375, 4700.22265625, 4672.39306640625, 4584.31982421875, 
    4010.41625976562, 3564.20483398438, 4735.14501953125, 5071.17041015625, 
    5071.17041015625, 5107.759765625, 5276.87939453125, 5213.1474609375, 
    4960.7373046875, 4196.50537109375, 4798.19384765625, 4996.40087890625, 
    4996.40087890625, 4976.4970703125, 5143.41858983545, 5170.2080078125, 
    5072.78857421875, 5198.359375, 5396.099609375, 5497.41015625, 5500, 5500, 
    5500, 5329.34130859375, 5473.99560546875, 5307.88232421875, 
    5297.4912109375, 5180.599609375, 5171.4072265625, 5293.05712890625, 
    5115.814453125, 5039.970703125, 5032.216796875, 4922.17333984375, 
    5124.61279296875, 4976.62451171875, 4852.5703125, 4794.8427734375, 
    4730.60595703125, 4709.47216796875, 4621.880859375, 4293.18310546875, 
    4116.666015625, 4153.27197265625, 4317.78125, 4198.8515625, 
    4293.060546875, 4293.060546875, 4357.39599609375, 4127.994140625, 
    4179.11669921875, 4008.75268554688, 3710.5302734375, 3570.740234375, 
    3362.02661132812, 3077.42333984375, 2832.45703125, 2692.38500976562, 
    2782.12329101562, 3108.04931640625, 3373.51733398438, 3516.03149414062, 
    3642.85668945312, 3864.67846679688, 3909.71728515625, 3937.41455078125, 
    4047.33178710938, 3958.9794921875, 3964.9990234375, 3964.9990234375, 
    3833.45434570312, 3709.1953125, 3644.75317382812, 3505.41552734375, 
    3168.72534179688, 3267.21630859375, 3078.98754882812, 3078.45874023438, 
    3270.23315429688, 3400.4970703125, 3519, 3664.58129882812, 
    3651.34521484375, 4000.61743164062, 4000.61743164062, 3925.3466796875, 
    4035.77880859375, 3960.64233398438, 4138.91259765625, 4129.89453125, 
    4136.90869140625, 4029.2314453125, 3990.11010742188, 3990.11010742188, 
    2946.39624023438, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 50, 80, 180, 1052.05932617188, 3579.77001953125, 
    4407.56787109375, 4973.09912109375, 5120.49267578125, 5212.51708984375, 
    5242.9677734375, 5203.673828125, 5176.759765625, 5167.44580078125, 
    5117.20556640625, 5115.03173828125, 5101.5615234375, 5088.56982421875, 
    5066.37548828125, 5012.69873046875, 5119.6015625, 5119.6015625, 
    4892.37353515625, 4962.9736328125, 4990.126953125, 4884.58349609375, 
    4669.59521484375, 4648.2255859375, 4548.634765625, 4270.94921875, 
    3729.97778320312, 3958.673828125, 4037.56030273438, 3772.69897460938, 
    3970.42919921875, 4004.35180664062, 4004.35180664062, 3997.69775390625, 
    3795.0361328125, 3553.30517578125, 3284.86083984375, 2764.11596679688, 
    2667.96923828125, 2714.431640625, 3015.197265625, 3165.44384765625, 
    3127.3291015625, 2985.67749023438, 3115.52978515625, 3311.52099609375, 
    3246.77612304688, 3182.03686523438, 3361.05859375, 3627.86010742188, 
    4102.2421875, 4341.826171875, 4585.45166015625, 4818.48681640625, 
    4937.98046875, 5121.3154296875, 5034.84716796875, 5034.84716796875, 
    5091.4921875, 5129.07666015625, 5111.65283203125, 5176.53076171875, 
    5248.443359375, 5216.47412109375, 5057.46728515625, 5063.58251953125, 
    5063.58251953125, 4685.55908203125, 4274.5966796875, 4419.18185522252, 
    4803.732421875, 4779.07571895829, 4818.68798828125, 4865.63134765625, 
    4852.9580078125, 5124.4912109375, 5097.3837890625, 5097.3837890625, 
    5009.75146484375, 4361.22021484375, 3555, 3555, 3215.22680664062, 
    3934.65405273438, 4225.9169921875, 4093.07592773438, 3946.86303710938, 
    3946.86303710938, 3746.876953125, 4794.759765625, 5488.634765625, 
    5347.3896484375, 4918.240234375, 4780.1826171875, 4644.82861328125, 
    4171.36474609375, 3994.51318359375, 3545.70654296875, 2454.45556640625, 
    2944.83276367188, 2997.72705078125, 2997.72705078125, 2045.44567871094, 
    2016.08728027344, 2548.26391601562, 3269.12646484375, 3163.03491210938, 
    3684.66723632812, 4270.1474609375, 4133.5869140625, 4603.2763671875, 
    4746.49072265625, 5235.111328125, 5256.1962890625, 5316.47509765625, 
    5293.291015625, 5292.00830078125, 5133.11328125, 4997.7890625, 
    4569.9150390625, 4537.16748046875, 4383.7021484375, 4297.7744140625, 
    4198.375, 4307.9609375, 4144.9658203125, 4324.396484375, 
    4273.38134765625, 4267.880859375, 4055.46655273438, 3688.6630859375, 
    2873.74975585938, 1287.97045898438, 2002.8291015625, 3177.78930664062,
  3330, 3639.09448242188, 3639.09448242188, 3585.81103515625, 3779.162109375, 
    3778.01245117188, 3781.765625, 3706.31372070312, 3578.6953125, 
    3794.52661132812, 3863.92822265625, 3836.57495117188, 3725.33349609375, 
    3852.3759765625, 4005.98413085938, 4106.0869140625, 4181.91015625, 
    4282.5146484375, 4375.7998046875, 4375.7998046875, 4492.27587890625, 
    4495.5185546875, 4687.6357421875, 4749.072265625, 4749.072265625, 
    4760.70947265625, 4760.70947265625, 4686.43212890625, 4856.21826171875, 
    4827.07763671875, 4738.73876953125, 4784.0615234375, 4784.0615234375, 
    4846.23193359375, 4896.2939453125, 5112.30810546875, 5039.064453125, 
    5118.01953125, 5095.93603515625, 5041.37255859375, 5261.373046875, 
    5256.0107421875, 5260.8994140625, 5444.48583984375, 5500, 5500, 
    5423.63818359375, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5494.71826171875, 5500, 5407.1552734375, 4689.56298828125, 
    1869.00341796875, 294.462890625, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    2671.00512695312, 4669.82568359375, 4763.9130859375, 4521.943359375, 
    4540, 4547.06201171875, 4490.27197265625, 4657.39111328125, 
    5027.3955078125, 4822.724609375, 4834.02099609375, 4823.8720703125, 
    3721.27612304688, 2341.13525390625, 1432.22448730469, 1616, 1616, 
    911.409484863281, 870.5537109375, 1186.11877441406, 1843.21069335938, 
    1792.85009765625, 1675.01892089844, 1009.32751464844, 150, -0, 200, 
    656.258728027344, 791.805480957031, 1870.53759765625, 3594.04907226562, 
    3594.04907226562, 4157.419921875, 5143.41858983545, 5457.27294921875, 
    5391.7041015625, 5327.82666015625, 5286.3857421875, 5143.41858983545, 
    5090.689453125, 4044.01904296875, 4458.166015625, 4458.166015625, 
    4735.14501953125, 5071.17041015625, 5387.13037109375, 5257.064453125, 
    5266.63134765625, 5213.974609375, 4891.50732421875, 4940.30615234375, 
    5297.71875, 5375.546875, 5409.52783203125, 5387.65673828125, 
    5377.8076171875, 5416.98486328125, 5242.662109375, 5422.7763671875, 5500, 
    5500, 5492.92822265625, 5397.51513671875, 5500, 5500, 5464.94091796875, 
    5173.583984375, 5088.42333984375, 5307.47314453125, 5178.22412109375, 
    5143.41858983545, 5034.1708984375, 4955.42919921875, 4866.1025390625, 
    4808.75390625, 4891.69677734375, 4779.07571895829, 4728.0166015625, 
    4547.67431640625, 4539.1650390625, 4463.05224609375, 4372.6103515625, 
    4177.71728515625, 4051.001953125, 4315.3544921875, 4339.35595703125, 
    3903.14306640625, 4293.060546875, 4293.060546875, 3614.8935546875, 
    4034.41772460938, 4034.41772460938, 4006.1435546875, 3710.5302734375, 
    3245.615234375, 2856.85400390625, 2857.74682617188, 2558.36376953125, 
    2482.87841796875, 2705.419921875, 3107.73901367188, 3413.16162109375, 
    3507.544921875, 3629.1865234375, 3815.43383789062, 3866.68481445312, 
    4002.13671875, 3727.85546875, 3635.10083007812, 3561.39038085938, 
    3623.59375, 3587.1650390625, 3389.79345703125, 3306.25952148438, 
    3192.96557617188, 2918.59936523438, 3076.24145507812, 3329.78588867188, 
    3455.81274414062, 3577.06567382812, 3502.45336914062, 3781.34790039062, 
    3968.68383789062, 3678.54638671875, 3988.73266601562, 3988.73266601562, 
    3872.69458007812, 3867.23461914062, 3987.25537109375, 3959.419921875, 
    4001.90258789062, 4029.2314453125, 4036.39526367188, 3990.11010742188, 
    3990.11010742188, 3872.95190429688, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 40, 90, 685.862060546875, 
    2398.02319335938, 3758.19653320312, 4292.69091796875, 4757.27685546875, 
    5031.96875, 5090.845703125, 5115.94140625, 5124.4130859375, 
    5124.4130859375, 5089.24658203125, 5051.6865234375, 5045.58349609375, 
    5038.2099609375, 5018.22216796875, 4996.78369140625, 4886.3583984375, 
    4874.9169921875, 4861.2890625, 4934.3388671875, 4761.6845703125, 
    4650.30126953125, 4621.3466796875, 4450.9912109375, 4150, 
    4012.36401367188, 4012.36401367188, 4304.58251953125, 4193.6640625, 
    4180.4111328125, 4106.91552734375, 4020.27392578125, 4004.35180664062, 
    3837.8505859375, 3832.56420898438, 3694.3818359375, 3291.11010742188, 
    2900.69750976562, 2878.02783203125, 3101.00830078125, 3325.06225585938, 
    3325.06225585938, 2175.15209960938, 3512.63427734375, 3512.63427734375, 
    3249.5068359375, 3155.59716796875, 3193.55102539062, 3361.05859375, 
    3627.86010742188, 3721.27612304688, 3876.33032226562, 3127.033203125, 
    4808.2265625, 4971.68896484375, 4999.2568359375, 5039.0703125, 
    5034.84716796875, 5032.5009765625, 5028.2197265625, 5009.81982421875, 
    4906.9306640625, 4993.20751953125, 4959.80615234375, 5057.46728515625, 
    5063.58251953125, 5063.58251953125, 5087.71826171875, 4955.8515625, 
    4764.01416015625, 4712.59765625, 4578.53857421875, 4487.7265625, 
    4603.46044921875, 4065.89147763595, 4046.32006835938, 4290.22509765625, 
    4317.28173828125, 4361.22021484375, 4361.22021484375, 3555, 3555, 
    3256.833984375, 3832.24682617188, 4419.18185522252, 4426.83447265625, 
    4185.68505859375, 4184.2724609375, 3803.17407226562, 4120.85888671875, 
    5143.759765625, 5467.18505859375, 5227.68017578125, 5157.673828125, 
    4890.22021484375, 4626.66455078125, 4459.66943359375, 4080.26171875, 
    2901.2412109375, 2944.83276367188, 3161.06518554688, 3277.81909179688, 
    3277.81909179688, 2706.87109375, 2350.83422851562, 1947.86096191406, 
    2650.98583984375, 3198.912109375, 3656.25830078125, 3865.06201171875, 
    4479.4501953125, 4756.38916015625, 5157.08935546875, 5168.5966796875, 
    5161.03076171875, 5159.11865234375, 5170.3779296875, 5049.255859375, 
    4872.89599609375, 4568.01904296875, 4368.828125, 4338.4326171875, 
    4275.287109375, 4170.69580078125, 4204.28076171875, 4319.0009765625, 
    4385.412109375, 4188.3037109375, 4190.48681640625, 3976.50415039062, 
    3688.6630859375, 3309.67724609375, 2645.9970703125, 1711.14599609375, 
    2054.68505859375,
  2353.56079101562, 3639.09448242188, 3903.4970703125, 3874.19384765625, 
    3911.05004882812, 3984.81665039062, 3898.85522460938, 3870.98852539062, 
    3832.46142578125, 3849.3671875, 4015.89892578125, 4054.39135742188, 
    3885.57739257812, 4032.0205078125, 4273.72705078125, 4099.83447265625, 
    4373.42724609375, 4427.2392578125, 4477.2666015625, 4375.7998046875, 
    4517.4189453125, 4674.87646484375, 4687.6357421875, 4826.94921875, 
    4949.63037109375, 4760.70947265625, 4971.080078125, 5053.42529296875, 
    5053.42529296875, 4817.0185546875, 4919.4501953125, 4948.9794921875, 
    5109.5947265625, 5109.5947265625, 5100.31201171875, 5077.45068359375, 
    4946.689453125, 4756.1748046875, 4804.61474609375, 5041.37255859375, 
    5207.046875, 5347.46875, 5310.72216796875, 5416.34912109375, 
    5407.19921875, 5486.16455078125, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5189.37109375, 5029.751953125, 4004.232421875, 931.482116699219, 
    70, 50, 50, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 2273.92333984375, 
    4669.82568359375, 4749.64013671875, 4659.2119140625, 4540, 
    4661.30615234375, 4103.498046875, 4593.04248046875, 4791.33935546875, 
    4975.81689453125, 4481.9716796875, 3545.7861328125, 2842.02685546875, 
    2341.13525390625, 1373.11779785156, 1616, 1616, 1760.74377441406, 
    1760.74377441406, 1616.94702148438, 1792.85009765625, 1851.72729492188, 
    1635.947265625, 1009.32751464844, -0, 40, 1336.12280273438, 2380, 
    2417.80834960938, 2385.90893554688, 4395.34619140625, 4631.61083984375, 
    5500, 5500, 5500, 5500, 5460.79833984375, 5291.26904296875, 
    5185.75439453125, 5090.689453125, 4679.7626953125, 4700.81005859375, 
    4700.81005859375, 4278.0380859375, 5052.77587890625, 5390.90966796875, 
    5293.734375, 5317.84375, 5237.11572265625, 5160.4541015625, 
    5117.3623046875, 5226.44384765625, 5386.6279296875, 5500, 
    5444.25927734375, 5444.369140625, 5500, 5486.0185546875, 5500, 5500, 
    5369.58642578125, 5319.47509765625, 5300.62646484375, 5386.85400390625, 
    5421.64111328125, 5235.92578125, 5101.60302734375, 5088.42333984375, 
    5033.28271484375, 4898.25, 4913.390625, 4883.95068359375, 
    4738.44384765625, 4666.5654296875, 4730.50146484375, 4716.7978515625, 
    4543.79052734375, 4566.923828125, 4373.65673828125, 4378.99169921875, 
    4284.1328125, 4311.98583984375, 4115.86767578125, 3924.51782226562, 
    3919.98046875, 3938.5244140625, 3991.7431640625, 4082.8779296875, 
    4295.63671875, 3788.9658203125, 3901.93359375, 3901.93359375, 
    3945.83813476562, 3565.70288085938, 3206.48510742188, 2719.9873046875, 
    2758.41088867188, 2804.79443359375, 2904.32641601562, 2778.70288085938, 
    3160.38354492188, 3446.302734375, 3517.14331054688, 3598.423828125, 
    3606.13842773438, 3678.56616210938, 3494.4638671875, 3306.1865234375, 
    3135.82177734375, 3283.46606445312, 3522.55078125, 3599.46362304688, 
    3207.0087890625, 3281.21411132812, 3008.10375976562, 3247.00146484375, 
    3362.08349609375, 3366.85131835938, 3653.40795898438, 3600.70141601562, 
    3727.44091796875, 3907.1044921875, 3953.30541992188, 3678.54638671875, 
    3700.400390625, 3968.06518554688, 3880.41796875, 3868.4892578125, 
    3970.51171875, 4046.93823242188, 4038.97973632812, 3994.00439453125, 
    3994.00439453125, 3979.9404296875, 4065.89147763595, 4065.89147763595, 
    425.785466617812, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 40, 40, 80, 770.675598144531, 2723.22119140625, 3721.27612304688, 
    4339.283203125, 4670.103515625, 4794.4072265625, 4933.27734375, 
    4998.26220703125, 5019.45703125, 4974.4775390625, 4967.87158203125, 
    4972.48583984375, 4961.67431640625, 4933.7509765625, 4970.12255859375, 
    4995.46240234375, 4928.81103515625, 4828.1787109375, 4813.2119140625, 
    4500.083984375, 4586.017578125, 4353.0205078125, 4307.52490234375, 
    4358.8154296875, 4366.1162109375, 4370.53271484375, 4301.1962890625, 
    4314.16455078125, 4159.3720703125, 4156.5537109375, 3881.7353515625, 
    3850.71264648438, 3940.93408203125, 3900.63061523438, 3526.24609375, 
    2914.45385742188, 2700.9501953125, 3002.43383789062, 3273.806640625, 
    3444.36547851562, 3523.62841796875, 3682.91381835938, 3682.91381835938, 
    3680.48217773438, 3680.48217773438, 3633.2275390625, 3193.55102539062, 
    3361.05859375, 3627.86010742188, 4015.0947265625, 4252.62353515625, 
    4402.83056640625, 4763.14501953125, 5002.580078125, 5072.791015625, 
    5120.546875, 5034.84716796875, 5222.75732421875, 5190.22021484375, 
    5118.36572265625, 4991.64111328125, 4653.748046875, 4987.0009765625, 
    5013.2275390625, 5063.58251953125, 5064.36865234375, 4975.4921875, 
    4889.17529296875, 4764.01416015625, 4760.2470703125, 4483.17578125, 
    4252.5341796875, 3867.91845703125, 2858.5751953125, 270.610395222517, 
    326.990295410156, 2211.01147460938, 3290.22924804688, 3290.22924804688, 
    3582.31616210938, 3582.31616210938, 4374.2724609375, 4710.38623046875, 
    4712.69873046875, 4590.5625, 4274.12939453125, 4134.95751953125, 
    3766.7333984375, 3567.71264648438, 5045.86181640625, 5500, 
    5390.0048828125, 5168.923828125, 5046.4697265625, 4852.3076171875, 
    4851.1298828125, 4365.4208984375, 3304.15112304688, 2434.76806640625, 
    3161.06518554688, 3648.7734375, 3697.50048828125, 3687.35424804688, 
    3452.61254882812, 3250.61181640625, 3224.99536132812, 3492.28271484375, 
    3656.25830078125, 3792.30737304688, 4089.12109375, 4450.2587890625, 
    4539.330078125, 5062.58203125, 4959.857421875, 4959.857421875, 
    4958.52978515625, 4715.97119140625, 4520.6708984375, 4453.32666015625, 
    4315.6728515625, 4270.3876953125, 4305.1669921875, 4351.11181640625, 
    4330.6220703125, 4353.68896484375, 4361.4189453125, 4207.810546875, 
    4069.205078125, 3957.11645507812, 3643.50390625, 3321.02612304688, 
    2969.36352539062, 2564.14819335938, 2492.04321289062,
  2902.29736328125, 3016.46337890625, 3721.27612304688, 3825.22094726562, 
    4003.35400390625, 3895.14233398438, 3981.2314453125, 3895.947265625, 
    3988.94921875, 3970.83935546875, 3851.00439453125, 3915.53564453125, 
    4046.69360351562, 4195.46533203125, 4436.671875, 4484.0732421875, 
    4541.28125, 4618.27587890625, 4572.43896484375, 4375.7998046875, 
    4522.82568359375, 4673.14794921875, 4552.40771484375, 5004.96435546875, 
    5004.96435546875, 5004.96435546875, 4874.8359375, 5233.24609375, 
    5434.04833984375, 4817.0185546875, 4894.283203125, 4948.9794921875, 
    5109.5947265625, 5109.5947265625, 4508.1513671875, 3399.8466796875, 
    1877.72021484375, 1224.30883789062, 2295.63720703125, 4248.2626953125, 
    4673.01708984375, 4673.01708984375, 4664.90087890625, 4748.78173828125, 
    4812.77587890625, 4953.681640625, 5219.7666015625, 5181.3212890625, 
    5233.3251953125, 5119.2265625, 4649.29296875, 3126.49780273438, 
    2005.56457519531, 1697.12502302956, 1746.70434570312, 230, 90, 0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 100, 4439.56787109375, 
    4815.31494140625, 4877.73193359375, 4513.5478515625, 4610, 
    4612.96630859375, 4650.57470703125, 4694.58740234375, 4694.58740234375, 
    3131.73510742188, 2861.56469726562, 2337.43359375, 1572.04309082031, 
    1059.37036132812, 1616, 1833.28149414062, 1833.28149414062, 
    1760.74377441406, 1616.94702148438, 1589.40393066406, 1589.40393066406, 
    765.529602050781, -0, -0, 586.903503417969, 2177.28369140625, 2380, 
    2385.90893554688, 2385.90893554688, 4395.34619140625, 5500, 5500, 5500, 
    5445.0703125, 5500, 5425.6201171875, 5296.29248046875, 4857.06298828125, 
    3687.05883789062, 4966.00927734375, 5005.8681640625, 5059.8759765625, 
    5094.2919921875, 5128.048828125, 5322.38623046875, 5382.1337890625, 
    5389.13818359375, 5392.04248046875, 5273.94287109375, 5117.3623046875, 
    5279.5107421875, 5329.95361328125, 5338.58154296875, 5435.19140625, 
    5483.8134765625, 5442.9521484375, 5416.65283203125, 5493.01171875, 
    5226.1015625, 4995.10546875, 4969.421875, 5009.17138671875, 
    5009.17138671875, 5131.23291015625, 5115.61376953125, 5101.60302734375, 
    5047.08935546875, 4633.779296875, 4743.24560546875, 4756.767578125, 
    4756.767578125, 4601.6103515625, 4611.16796875, 4673.01318359375, 
    4451.38525390625, 4286.3037109375, 4104.8779296875, 4044.6435546875, 
    4017.34228515625, 4036.13940429688, 4046.20678710938, 3811.26318359375, 
    3819.34594726562, 3949.4384765625, 4005.0224609375, 3992.86767578125, 
    4169.8125, 4217.82861328125, 3788.9658203125, 3543.41015625, 
    3319.4931640625, 2951.39086914062, 3328.2978515625, 3328.2978515625, 
    3205.45532226562, 3029.0947265625, 2804.79443359375, 2983.86254882812, 
    2841.04028320312, 3094.90209960938, 3481.30639648438, 3387.2978515625, 
    3488.99780273438, 3395.00024414062, 3477.69848632812, 3146.05688476562, 
    3078.73022460938, 3183.15014648438, 3327.33959960938, 3660.54296875, 
    3650.90747070312, 3527.85083007812, 3387.2978515625, 3397.71459960938, 
    3415.55004882812, 3293.86694335938, 3424.34106445312, 3644.41357421875, 
    3600.70141601562, 3887.37084960938, 3962.98193359375, 4003.05029296875, 
    4052.3525390625, 3948.35229492188, 3961.89331054688, 3893.18090820312, 
    3819.23193359375, 3974.275390625, 3947.27392578125, 3981.99487304688, 
    4038.33227539062, 4005.1435546875, 4026.86938476562, 4161.8095703125, 
    4076.65502929688, 2544.74365234375, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 40, 40, 40, 70, 733.100463867188, 
    2656.07983398438, 3641.06640625, 4295.40576171875, 4652.3544921875, 
    4803.30908203125, 4861.794921875, 4835.61474609375, 4871.96923828125, 
    4898.6572265625, 4888.1845703125, 4845.18603515625, 4791.22412109375, 
    4856.6083984375, 4882.4443359375, 4758.9892578125, 4606.6201171875, 
    4657.14892578125, 4455.373046875, 4459.111328125, 4353.0205078125, 
    4140.27734375, 4171.49462890625, 4394.27392578125, 4366.1162109375, 
    4249.716796875, 4087.04370117188, 4040.96948242188, 4021.14086914062, 
    3916.2333984375, 3683.48950195312, 3694.2578125, 3694.2578125, 
    3543.8662109375, 3414.03442382812, 2986.38549804688, 3002.43383789062, 
    3315.26000976562, 3477.07348632812, 3711.24731445312, 3682.91381835938, 
    3800.9052734375, 3840.14477539062, 3834.4267578125, 3943.22412109375, 
    3867.7607421875, 3984.6103515625, 3242.10522460938, 3509.56298828125, 
    4090.3359375, 4402.83056640625, 4630.15283203125, 4704.61181640625, 
    4848.80615234375, 4854.1064453125, 5007.78271484375, 5277.6796875, 
    5279.74560546875, 5231.15087890625, 5221.82861328125, 5097.4208984375, 
    5053.07421875, 5079.7978515625, 5044.427734375, 5021.89306640625, 
    4884.21923828125, 4498.916015625, 4675.64501953125, 4675.64501953125, 
    4124.14208984375, 3366.96337890625, 1989.63879394531, 210, 210, 210, 
    397.158264160156, 1681.00024414062, 2410.22094726562, 3582.31616210938, 
    3582.31616210938, 4374.2724609375, 4503.38623046875, 4492.1396484375, 
    4587.81396484375, 4274.12939453125, 3926.86767578125, 3817.41137695312, 
    3558.06079101562, 3721.27612304688, 5463.20556640625, 5413.68505859375, 
    5319.7373046875, 5328.66650390625, 5034.06298828125, 4878.28369140625, 
    4365.4208984375, 3304.15112304688, 2434.76806640625, 3178.15966796875, 
    3463.7705078125, 3721.27612304688, 3880.67724609375, 3682.2734375, 
    3873.06323242188, 3867.77954101562, 3867.77954101562, 3492.28271484375, 
    3068.4755859375, 3810.3427734375, 4127.0869140625, 4408.47265625, 
    4868.92578125, 4993.7578125, 4914.796875, 5026.6171875, 4642.57373046875, 
    4387.66943359375, 4348.91455078125, 4407.50341796875, 4292.150390625, 
    4376.0576171875, 4246.84716796875, 4330.6220703125, 4345.92822265625, 
    4220.71044921875, 4159.107421875, 4086.36962890625, 3826.26831054688, 
    3640.63720703125, 3286.72241210938, 2969.36352539062, 2863.84448242188, 
    2910,
  2910, 2912.04223632812, 3012.11376953125, 3402.01513671875, 
    3810.38403320312, 3822.76806640625, 3387.537109375, 3700.95434570312, 
    4026.1572265625, 4047.8505859375, 4022.77954101562, 4219.6845703125, 
    4315.54296875, 4345.88232421875, 4419.18185522252, 4497.58935546875, 
    4515.2431640625, 4579.3427734375, 4512.03857421875, 4296.583984375, 
    4419.18185522252, 4419.18185522252, 4572.626953125, 5273.59765625, 5500, 
    5500, 5282.8154296875, 5249.5068359375, 5224.46630859375, 
    4545.5009765625, 2405, 2715, 2719.88940429688, 2719.88940429688, 
    536.623229980469, 40, -0, -0, -0, 120, 629.9306640625, 629.9306640625, 
    270.610395222517, 284.156616210938, 2889.74853515625, 3857.99658203125, 
    3954.35717773438, 3954.35717773438, 3961.4228515625, 3428.0673828125, 
    1649.4208984375, 1342.57861328125, 845.124450683594, 110, 100, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 1680.57434082031, 
    4881.45263671875, 4881.86572265625, 4808.7685546875, 4719.919921875, 
    4691.974609375, 4638.77197265625, 4675.37109375, 4348.51904296875, 
    2384.02563476562, 2193.50732421875, 1133.11474609375, 1186.46875, 2535, 
    2533.82641601562, 2533.82641601562, 1833.28149414062, 1697.12502302956, 
    1718.38391113281, 1667.48327636719, 1159.55200195312, 80, 
    763.756103515625, 1205.72924804688, 1726.31384277344, 2296.76416015625, 
    2649.35375976562, 2649.35375976562, 1790.76647949219, 3699.3037109375, 
    5500, 5500, 5500, 5500, 5500, 5500, 5337.939453125, 4857.06298828125, 
    4811.57958984375, 5295.521484375, 5223.8505859375, 5180.6982421875, 
    5285.45751953125, 5128.048828125, 5425.90380859375, 5408.49560546875, 
    5498.28369140625, 5321.71044921875, 5181.7314453125, 5223.59423828125, 
    5285.81298828125, 5399.87060546875, 5305.2099609375, 5264.798828125, 
    5243.9619140625, 5300.71533203125, 5389.51025390625, 5295.3564453125, 
    5220.5283203125, 5148.44775390625, 5013.82958984375, 5250.01953125, 
    5144.5224609375, 5009.1845703125, 5063.26171875, 5063.26171875, 
    4785.47900390625, 4960.1943359375, 4877.13427734375, 4756.767578125, 
    4756.767578125, 4672.02294921875, 4593.87646484375, 4502.95458984375, 
    4465.80126953125, 4216.00146484375, 4119.162109375, 3090.14111328125, 
    3089.53784179688, 3198.2060546875, 3696.73803710938, 3696.73803710938, 
    3501.64990234375, 3621.49853515625, 3980.93725585938, 3969.8544921875, 
    3850.93896484375, 3190.048828125, 3543.41015625, 3629.169921875, 
    3629.169921875, 3623.51806640625, 3328.2978515625, 3328.2978515625, 
    3205.45532226562, 3029.0947265625, 2678.96752929688, 2867.72485351562, 
    3035.35034179688, 2927.83618164062, 3044.19970703125, 3246.07446289062, 
    3255.91259765625, 3343.4697265625, 3298.72216796875, 3327.16845703125, 
    3287.94848632812, 3287.94848632812, 3507.50659179688, 3566.9541015625, 
    3571.32446289062, 3496.59326171875, 3462.77758789062, 3392.19140625, 
    3593.9169921875, 3574.30029296875, 3587.96533203125, 3587.96533203125, 
    3645.42578125, 3842.74438476562, 3904.62133789062, 3928.4287109375, 
    3901.26098632812, 4001.40063476562, 3943.54321289062, 3859.25463867188, 
    3828.349609375, 3722.15454101562, 3813.1015625, 3972.4892578125, 
    3991.24926757812, 4005.1435546875, 4035.15161132812, 4076.65502929688, 
    4104.69384765625, 3908.916015625, 1252.89831542969, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 0, -0, -0, -0, -0, 40, 80, 
    1352.37316894531, 2873.84594726562, 3473.0322265625, 4030.47265625, 
    4531.03076171875, 4669.8974609375, 4765.96240234375, 4758.8076171875, 
    4722.27197265625, 4681.64208984375, 4676.45556640625, 4713.56640625, 
    4757.87060546875, 4757.87060546875, 4596.70947265625, 4701.765625, 
    4409.021484375, 4443.7763671875, 4474.7548828125, 4310.294921875, 
    3745.71704101562, 2855.03149414062, 4146.94677734375, 4249.716796875, 
    4355.25537109375, 4150, 3922.14379882812, 3980.57348632812, 
    3941.56420898438, 3883.56127929688, 3762.68237304688, 3760.04272460938, 
    3634.49487304688, 3514.3193359375, 3481.2744140625, 3281.19067382812, 
    2715.2294921875, 2991.193359375, 3321.546875, 3627.1494140625, 
    3883.61303710938, 4029.42944335938, 4104.41943359375, 4144.0234375, 
    3913.81787109375, 3913.81787109375, 3808.63793945312, 3304.4765625, 
    2768.744140625, 4046.17163085938, 3988.42016601562, 3988.42016601562, 
    3945.318359375, 4871.0947265625, 4911.7919921875, 5019.75732421875, 
    5217.7265625, 5236.6552734375, 5292.662109375, 5196.03076171875, 
    5082.55859375, 5044.427734375, 5054.93798828125, 4892.9501953125, 
    4794.14111328125, 4638.58984375, 4543.58154296875, 4399.056640625, 
    3694.48022460938, 1771.95861816406, 170, 130, 130, 130, 130, 130, 130, 
    664.643737792969, 2173.755859375, 3784.3193359375, 4065.89147763595, 
    4216.07763671875, 4161.2841796875, 4195.455078125, 2706.17431640625, 
    2600, 2640.5673828125, 2802.65576171875, 4903.63623046875, 
    5387.4130859375, 5269.25, 5267.3447265625, 5034.06298828125, 
    5045.80615234375, 4365.4208984375, 2288.26806640625, 1592.96484375, 
    1635.28515625, 2540.75854492188, 3742.4541015625, 3987.97729492188, 
    4080.22631835938, 4105.50146484375, 4105.50146484375, 4100.28662109375, 
    3506.34985351562, 2900.83618164062, 3170.63256835938, 3466.30810546875, 
    4267.7841796875, 4085.27099609375, 4720.3271484375, 5025.40185546875, 
    4839.9384765625, 4696.27587890625, 4547.93896484375, 4515.40673828125, 
    4666.5, 4510.85498046875, 4635.56494140625, 4513.62841796875, 
    4363.62451171875, 4324.0517578125, 4343.6650390625, 4220.8701171875, 
    4215.37353515625, 3867.65795898438, 3554.94897460938, 3286.72241210938, 
    2908.3681640625, 2773.57543945312, 2912.3876953125,
  3475.32641601562, 3466.5966796875, 3043.54443359375, 3597.32104492188, 
    3454.27465820312, 3620.46533203125, 3092.37231445312, 2910.86791992188, 
    3549.30981445312, 3887.25561523438, 4022.77954101562, 4279.724609375, 
    4347.001953125, 4345.88232421875, 4459.77734375, 4437.02587890625, 
    4316.50927734375, 4294.27001953125, 4296.583984375, 4296.583984375, 
    4500.38427734375, 4419.18185522252, 4572.626953125, 5361.61767578125, 
    5243.2373046875, 5440.9912109375, 5331.48828125, 4981.955078125, 
    4981.955078125, 3853.87670898438, 2414.18701171875, 2930.51586914062, 
    2925.40112304688, 2843.58984375, 476.123931884766, 40, -0, -0, -0, -0, 
    -0, -0, -0, -0, 60, 120, 718.495483398438, 698.805969238281, 
    698.805969238281, 536.538879394531, 536.538879394531, 336.698089599609, 
    120, 110, 60, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 50, 3224.55224609375, 4862.99365234375, 4822.0595703125, 
    4852.25537109375, 4544.05908203125, 4258.19482421875, 3291.05322265625, 
    3288.74658203125, 1847.90930175781, 1540.79467773438, 712.393676757812, 
    942.839303029559, 2883.76318359375, 2883.76318359375, 2533.82641601562, 
    1640.66259765625, 1983.26416015625, 1962.50537109375, 1711.50915527344, 
    1711.50915527344, 1670, 2046.23217773438, 2703.99096679688, 
    2996.44116210938, 2918.509765625, 3015.73461914062, 2674.5302734375, 
    2349.88818359375, 2287.62866210938, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 3758.16674804688, 5393.70556640625, 5272.46630859375, 
    5439.857421875, 5344.62744140625, 5289.8291015625, 5500, 
    5351.89501953125, 5500, 5486.78173828125, 5148.1416015625, 
    5144.01318359375, 5257.83154296875, 5288.5654296875, 5469.7509765625, 
    5369.17626953125, 5300.4921875, 5170.51123046875, 5218.29248046875, 
    5167.607421875, 5201.55322265625, 5308.75830078125, 5253.5498046875, 
    5013.82958984375, 5146.60205078125, 5143.41858983545, 5100.94287109375, 
    5115.96337890625, 5115.96337890625, 5072.11181640625, 4865.8701171875, 
    4881.1640625, 4726.2548828125, 4740.81884765625, 4672.02294921875, 
    4560.0341796875, 4627.84423828125, 4574.9052734375, 4393.611328125, 
    4193.75244140625, 3869.02075195312, 3560.19091796875, 3545.04541015625, 
    3658.99047851562, 3658.99047851562, 3501.64990234375, 3621.49853515625, 
    3660.58349609375, 3660.58349609375, 3658.63525390625, 3190.048828125, 
    3490.2841796875, 3656.41772460938, 3629.169921875, 3623.51806640625, 
    3094.259765625, 3196.31030273438, 2770.71020507812, 2833.17822265625, 
    2623.83618164062, 2902.86157226562, 2916.04931640625, 2917.91333007812, 
    3188.00854492188, 3137.9736328125, 3138.8232421875, 3270.73461914062, 
    2983.0634765625, 3194.16186523438, 3486.572265625, 3520.98876953125, 
    3621.9638671875, 3586.31127929688, 3592.60571289062, 3514.99780273438, 
    3667.51123046875, 3699.0263671875, 3699.0263671875, 3674.7041015625, 
    3674.07666015625, 3587.96533203125, 3660.21850585938, 3724.72143554688, 
    3744.79418945312, 3943.12231445312, 3788.12036132812, 3926.80517578125, 
    3955.63720703125, 3868.13745117188, 3967.01489257812, 3849.93432617188, 
    3389.6640625, 3463.45581054688, 2447.24584960938, 2427.92846679688, 
    4129.3740234375, 4236.08740234375, 3908.916015625, 3908.916015625, 
    2802.548828125, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 40, 230, 962.111145019531, 2303.4638671875, 
    3189.99584960938, 3624.3515625, 3884.95727539062, 4043.302734375, 
    4200.48486328125, 4318.0205078125, 4491.2919921875, 4589.185546875, 
    4663.51171875, 4689.78076171875, 4493.3681640625, 4562.42724609375, 
    4447.85791015625, 4285.51904296875, 4305.0693359375, 4279.9609375, 
    3734.93383789062, 3604.630859375, 2408.87524414062, 4150, 
    4065.89147763595, 4304.44921875, 4308.24462890625, 4264.09375, 
    4309.22216796875, 4302.50537109375, 4071.2255859375, 3877.53784179688, 
    3731.8779296875, 3721.40991210938, 3581.82836914062, 3399.78295898438, 
    3281.19067382812, 3276.44873046875, 3097.82397460938, 3280.71533203125, 
    3557.92333984375, 3797.02880859375, 4029.42944335938, 4105.00439453125, 
    4191.5693359375, 3913.81787109375, 3952.93530273438, 4018.32861328125, 
    3483.89575195312, 2853.083984375, 2892.8447265625, 2892.8447265625, 
    2669.7587890625, 3945.318359375, 4079.63232421875, 4079.63232421875, 
    4950.4755859375, 5017.12841796875, 5218.43359375, 5228.056640625, 
    5207.70947265625, 5082.55859375, 5021.67333984375, 4941.95556640625, 
    4724.5107421875, 4543.07666015625, 4313.34228515625, 4142.28955078125, 
    3730.041015625, 2225.87084960938, 443.4267578125, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 404.1171875, 3013.77368164062, 3677.96411132812, 
    3811.099609375, 3906.77197265625, 3609.01904296875, 2334.91650390625, 
    2250, 2250, 4153.466796875, 5126.29833984375, 5126.29833984375, 
    5131.9873046875, 5013.4111328125, 5003.3095703125, 4163.703125, 
    1554.60375976562, 899.838500976562, 1284.9208984375, 2638.43310546875, 
    3606.97143554688, 4000.63842773438, 4206.48193359375, 4310.6826171875, 
    4283.96435546875, 4283.96435546875, 4251.912109375, 3652.82299804688, 
    2945.76416015625, 3044.37255859375, 4003.38793945312, 4189.30859375, 
    4720.3271484375, 4870.00830078125, 5049.15234375, 4682.41162109375, 
    4707.2822265625, 4759.67236328125, 4679.306640625, 4622.59423828125, 
    4670.5458984375, 4511.083984375, 4507.70263671875, 4368.71826171875, 
    4324.0517578125, 4073.1669921875, 3991.64379882812, 3806.08984375, 
    3370.09497070312, 3200.57495117188, 2908.3681640625, 3049.21508789062, 
    3144.45385742188,
  3625.96362304688, 3543.5673828125, 2725.625, 2881.39965820312, 
    2881.39965820312, 2915.2080078125, 2915.2080078125, 2092.2900390625, 
    3312.91967773438, 3775.0732421875, 4022.77954101562, 4258.3828125, 
    4404.71923828125, 4340.39453125, 4340.39453125, 3865.935546875, 
    3865.935546875, 3189.7548828125, 3749.45190429688, 3923.93774414062, 
    3227.1884765625, 3349.95458984375, 4455.01416015625, 5350.13525390625, 
    5378.6298828125, 4764.6650390625, 4945.3173828125, 5336.62744140625, 
    5413.67822265625, 5182.287109375, 4779.07571895829, 4905.181640625, 
    4639.6474609375, 4294.17236328125, 1232.86547851562, 40, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 50, 50, 50, 60, 60, 60, 40, 40, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 70, 
    4361.3505859375, 4803.70751953125, 4875.6240234375, 4072.728515625, 
    3090.29321289062, 3288.74658203125, 3343.15356445312, 1503.84399414062, 
    1418.45043945312, 944.09814453125, 1377.20825195312, 2883.76318359375, 
    2883.76318359375, 1034.09033203125, 962.455749511719, 1998.14489746094, 
    3654.84497070312, 3559.60571289062, 3046.75537109375, 1669.72204589844, 
    2527.96533203125, 3637.87768554688, 3686.42211914062, 3686.42211914062, 
    3582.0234375, 2349.88818359375, 2349.88818359375, 2405.54516601562, 
    3966.87329101562, 5500, 5500, 5478.0068359375, 5500, 5500, 5500, 
    4796.5751953125, 5467.35302734375, 5500, 5500, 5500, 5143.41858983545, 
    5220.5146484375, 5282.298828125, 5482.78857421875, 5349.37158203125, 
    5302.86572265625, 5500, 5383.3740234375, 5452.5888671875, 
    5443.5517578125, 5423.5634765625, 5230.7490234375, 5209.90283203125, 
    5166.19970703125, 5155.2373046875, 5031.2509765625, 5143.41858983545, 
    5171.22900390625, 4998.9306640625, 4674.6708984375, 5084.86865234375, 
    5100.94287109375, 5115.96337890625, 5128.7109375, 5062.54150390625, 
    4965.71484375, 4859.1552734375, 4726.2548828125, 4621.39013671875, 
    4450.29248046875, 4571.677734375, 4506.5947265625, 4356.57275390625, 
    4220.74853515625, 4240.5859375, 3869.02075195312, 3560.19091796875, 
    3600.44213867188, 3600.44213867188, 3189.462890625, 3617.927734375, 
    3500.68701171875, 3475.43627929688, 3489.65942382812, 3218.08911132812, 
    3089.103515625, 3281.79028320312, 3281.79028320312, 3482.08618164062, 
    3419.93359375, 3293.076171875, 3065.78548661781, 3034.39086914062, 
    2887.40991210938, 2661.41088867188, 2631.017578125, 2784.64624023438, 
    3026.52099609375, 3066.65112304688, 3240.68383789062, 3339.14038085938, 
    3376.03149414062, 3376.03149414062, 3595.92504882812, 3650.93408203125, 
    3666.96533203125, 3691.40161132812, 3804.24194335938, 3760.4814453125, 
    3653.16821289062, 3667.51123046875, 3770.67016601562, 3724.47900390625, 
    3246.453125, 3586.48828125, 3457.427734375, 3609.33666992188, 
    3456.60717773438, 3584.55883789062, 3785.95678710938, 3864.6279296875, 
    3936.47265625, 3862.62133789062, 3750.5068359375, 3855.67016601562, 
    3931.66528320312, 3959.09765625, 3951.06176757812, 4122.62109375, 
    4095.55834960938, 4183.4296875, 4252.8974609375, 3978.59252929688, 
    3789.29370117188, 3789.29370117188, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 60, 190, 1916.43872070312, 
    2952.29052734375, 3528.73364257812, 3857.21264648438, 4055.11401367188, 
    4043.302734375, 4042.85375976562, 4119.078125, 4322.80029296875, 
    4294.29052734375, 4294.29052734375, 4291.66162109375, 4291.66162109375, 
    3658.83081054688, 3087.96606445312, 3723.44482421875, 3852.955078125, 
    4046.49462890625, 3640.00219726562, 3640.00219726562, 4150, 4150, 
    4156.64013671875, 4358.146484375, 4264.09375, 4202.1826171875, 
    4381.619140625, 4094.845703125, 4054.15307617188, 3989.39208984375, 
    3741.53125, 3689.67041015625, 3528.525390625, 3469.31323242188, 
    3272.40698242188, 3184.80859375, 2895.88159179688, 3409.24145507812, 
    3546.65209960938, 3931.24536132812, 3963.255859375, 3963.255859375, 
    3959.9951171875, 3959.9951171875, 3952.93530273438, 4044.06787109375, 
    3999.3955078125, 3978.69311523438, 3666.58911132812, 2466.66776221529, 
    3668.40087890625, 3668.40087890625, 4291.4423828125, 4670.3466796875, 
    4883.98486328125, 5107.02001953125, 5107.02001953125, 4960.27978515625, 
    4932.39599609375, 4982.5546875, 4922.466796875, 4561.5263671875, 
    4078.7001953125, 3534.8896484375, 3373.26123046875, 2580.46948242188, 
    709.262573242188, 220, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    2660.65625, 3549.42993164062, 3634.5615234375, 3575.939453125, 
    3374.59643554688, 1913.32141113281, 1643.07507324219, 3426.3828125, 
    5092.052734375, 4996.953125, 5027.25146484375, 5018.50341796875, 
    4679.34912109375, 4083.22436523438, 1316.3330078125, 1174.67919921875, 
    1635.9150390625, 2855.53881835938, 3420.27587890625, 3682.0966796875, 
    3856.38330078125, 4122.23583984375, 4581.68017578125, 4745.86962890625, 
    4251.912109375, 4221.2861328125, 3923.56616210938, 4013.19409179688, 
    3452.84765625, 4276.6240234375, 4560.07470703125, 4618.37109375, 
    4618.37109375, 4725.65478515625, 4725.65478515625, 4725.65478515625, 
    4698.19091796875, 4680.66455078125, 4535.34423828125, 4516.65771484375, 
    4449.96240234375, 4387.45263671875, 4316.28271484375, 4166.78662109375, 
    3906.9228515625, 3744.927734375, 3370.09497070312, 3103.5263671875, 
    2814.08422851562, 3115.59692382812, 3613.73168945312,
  3981.9091796875, 3904.03344726562, 3791.23095703125, 3785.57861328125, 
    3785.57861328125, 3539.69995117188, 3018.76928710938, 1665.61022949219, 
    2141.47412109375, 3445.42846679688, 3961.89990234375, 4195.17236328125, 
    4334.630859375, 4243.74560546875, 2864.13110351562, 1390.68774414062, 
    2345.02954101562, 2345.02954101562, 2207.9921875, 2430.25659179688, 
    3193.5654296875, 3187.52172851562, 4733.29931640625, 5095.55712890625, 
    5095.55712890625, 4937.75146484375, 5079.77978515625, 5215.4453125, 
    5235.974609375, 5243.62255859375, 5144.31005859375, 5122.53173828125, 
    5080.841796875, 4863.81689453125, 1232.86547851562, 40, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    3034.5185546875, 4668.46630859375, 4668.46630859375, 4296.8037109375, 
    2814.6181640625, 2814.6181640625, 1724.60693359375, 1439.93896484375, 
    1174.64904785156, 1127.78625488281, 1377.20825195312, 2700, 2700, 
    1660.55432128906, 1939.81616210938, 2968.35229492188, 3559.60571289062, 
    3559.60571289062, 3046.75537109375, 1489.12023925781, 2585.2607421875, 
    3612.13134765625, 3705.20971679688, 4007.45166015625, 3978.93676757812, 
    3187.26000976562, 2350, 2350, 2350, 5500, 5500, 5496.07666015625, 5500, 
    5500, 4693.52099609375, 5500, 5500, 5500, 5500, 5428.70947265625, 
    5031.7685546875, 5066.94921875, 5066.94921875, 5335.625, 5407.021484375, 
    5315.05615234375, 5262.4228515625, 5173.443359375, 5335.7939453125, 
    5189.6689453125, 5332.7880859375, 5189.404296875, 5178.68994140625, 
    5102.13525390625, 5117.31396484375, 5036.4287109375, 5031.2509765625, 
    4704.12890625, 4704.12890625, 4751.240234375, 5009.1982421875, 
    4896.134765625, 4995.2421875, 5005.662109375, 4891.1669921875, 
    4815.58349609375, 4599.849609375, 4229.39013671875, 4131.9990234375, 
    4263.6494140625, 4305.5400390625, 4212.9140625, 4176.9208984375, 
    3906.0390625, 3906.0390625, 3837.79125976562, 3840.29125976562, 
    3658.1259765625, 3623.2919921875, 3873.88427734375, 3841.18041992188, 
    3898.10400390625, 3831.33837890625, 3570.76782226562, 3662.31762695312, 
    3534.41137695312, 3461.69409179688, 3469.76098632812, 3501.82763671875, 
    3500.35498046875, 3333.87036132812, 3239.13671875, 3034.39086914062, 
    2852.75366210938, 2727.35424804688, 2647.35034179688, 2821.32006835938, 
    3026.52099609375, 3094.05322265625, 3344.609375, 3369.64526367188, 
    3481.11254882812, 3683.16845703125, 3595.92504882812, 3650.93408203125, 
    3664.6953125, 3664.6953125, 3759.5234375, 3730.19702148438, 
    3653.16821289062, 3667.51123046875, 3803.5361328125, 3773.3046875, 
    3560.54028320312, 3480.76171875, 2995.62255859375, 2989.03881835938, 
    3441.271484375, 3780.07495117188, 3748.072265625, 3762.59033203125, 
    3970.6884765625, 3751.4072265625, 3891.75390625, 3888.45654296875, 
    3960.88208007812, 3931.8095703125, 4024.3798828125, 4124.17626953125, 
    4219.76708984375, 4094.3828125, 4215.78466796875, 4100.04736328125, 
    3966.21215820312, 3966.21215820312, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 90, 1351.30505371094, 
    2725.00854492188, 3185.64233398438, 3390.279296875, 3575.82421875, 
    3621.97827148438, 3640.20288085938, 4150, 4150, 4150, 4150, 
    3721.27612304688, 3258.4375, 2506.15966796875, 1579.4306640625, 
    1684.00329589844, 1895.50671386719, 2676.814453125, 3704.70288085938, 
    3704.70288085938, 4150, 4129.357421875, 4604.880859375, 4715.77734375, 
    4482.13916015625, 4419.18185522252, 4479.787109375, 4360.443359375, 
    4360.443359375, 4208.27587890625, 4027.44995117188, 3856.759765625, 
    3810.93896484375, 3637.43481445312, 3289.47509765625, 3131.49951171875, 
    2929.67626953125, 3145.25512695312, 3511.57568359375, 3768.87890625, 
    4035.71215820312, 3873.12719726562, 4034.06030273438, 4238.87841796875, 
    4385.2236328125, 4369.990234375, 3965.06762695312, 3965.06762695312, 
    3666.58911132812, 3553.45190429688, 3668.40087890625, 3668.40087890625, 
    2031.85363769531, 4670.3466796875, 4904.0966796875, 5107.02001953125, 
    5107.02001953125, 5031.84619140625, 4145.78857421875, 4908.38916015625, 
    4915.29833984375, 4378.169921875, 3876.05297851562, 3316.74780273438, 
    2762.26293945312, 1072.86096191406, 349.798828125, 160, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 2821.59448242188, 3161.12451171875, 
    3354.19702148438, 3339.51806640625, 2702.75048828125, 2250, 
    3550.18115234375, 5009.853515625, 4928.20263671875, 5017.41259765625, 
    4987.5986328125, 4722.29052734375, 3584.4169921875, 2006.02502441406, 
    2116.01904296875, 1935.05359591651, 2816.7998046875, 3420.27587890625, 
    4290.42431640625, 4583.81689453125, 4645.84814453125, 4682.51611328125, 
    4682.51611328125, 4238.15380859375, 4221.2861328125, 4390.302734375, 
    4390.302734375, 3368.4375, 3356.10107421875, 3505.53271484375, 4717.3125, 
    4618.37109375, 4725.65478515625, 4725.65478515625, 4725.65478515625, 
    4698.19091796875, 4543.2841796875, 4534.2802734375, 4487.69580078125, 
    4387.45263671875, 4387.45263671875, 4301.61767578125, 4052.2919921875, 
    3961.625, 3318.89721679688, 3249.17553710938, 3039.263671875, 
    3163.83447265625, 3252.60424804688, 3725.15258789062,
  3870.564453125, 3929.10498046875, 4006.07861328125, 4006.07861328125, 
    3807.63793945312, 3496.50146484375, 3258.71435546875, 2166.2275390625, 
    2077.07275390625, 1973.2333984375, 2262.49780273438, 2449.22387695312, 
    2154.32836914062, 2086.13818359375, 1806.37182617188, 2103.40576171875, 
    2731.37133789062, 2731.37133789062, 2207.9921875, 2711.27490234375, 
    3769.37451171875, 4395.07666015625, 4507.98583984375, 4743.6962890625, 
    4955.49951171875, 4917.25732421875, 5079.77978515625, 5122.6005859375, 
    5194.25341796875, 5361.1015625, 5298.11181640625, 5196.89697265625, 
    4995.56689453125, 4822.27978515625, 1003.23504638672, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 90, 
    4527.93896484375, 4720.9013671875, 4296.8037109375, 2692.88500976562, 
    2692.88500976562, 1941.92309570312, 1478.68884277344, 1312.4111328125, 
    1160.83044433594, 1337.00122070312, 2690.86279296875, 2766.02099609375, 
    2766.02099609375, 1939.81616210938, 2968.35229492188, 2969.9033203125, 
    2969.9033203125, 2376.04956054688, 1699.8759765625, 2585.2607421875, 
    3742.1962890625, 4169.0234375, 4236.51513671875, 3980.58984375, 
    3224.76000976562, 2098.17529296875, 2098.17529296875, 954.816955566406, 
    4390.9150390625, 5500, 5500, 5500, 5300.87451171875, 5500, 5500, 5500, 
    5500, 5407.74169921875, 5441.08251953125, 5449.99560546875, 
    5460.4638671875, 5212.8076171875, 5279.8330078125, 5202.2451171875, 
    5288.138671875, 5158.54345703125, 5192.82568359375, 5081.80615234375, 
    4925.798828125, 5003.7314453125, 5048.630859375, 5048.630859375, 
    5115.2353515625, 5096.083984375, 4985.42919921875, 4807.0380859375, 
    4515.0107421875, 4598.642578125, 4751.240234375, 4863.0068359375, 
    4865.6630859375, 4905.09423828125, 4846.3154296875, 4802.97314453125, 
    4419.18185522252, 4429.31689453125, 4124.74365234375, 4091.73388671875, 
    4042.916015625, 4175.9404296875, 4186.9755859375, 4073.09985351562, 
    4179.6884765625, 4282.2470703125, 4189.943359375, 4142.6884765625, 
    3926.8994140625, 3960.07446289062, 3942.68774414062, 3835.22509765625, 
    4011.1767578125, 3769.43872070312, 3794.65698242188, 3705.30419921875, 
    3684.4150390625, 3588.69970703125, 3534.84838867188, 3464.08276367188, 
    3449.92822265625, 3333.87036132812, 3262.75048828125, 2945.89526367188, 
    2946.18383789062, 2810.33276367188, 2697.96264648438, 2985.072265625, 
    3045.62426757812, 3196.9453125, 3200.92114257812, 3369.64526367188, 
    3523.63500976562, 3579.50561523438, 3489.63647460938, 3519.15942382812, 
    3564.50903320312, 3602.81372070312, 3611.49682617188, 3563.35302734375, 
    3600.36059570312, 3540.12377929688, 3690.3994140625, 3690.3994140625, 
    3704.1064453125, 3533.6240234375, 3297.63745117188, 3202.73413085938, 
    3706.076171875, 3761.04248046875, 3721.27612304688, 3763.1572265625, 
    3777.04296875, 3863.365234375, 3845.00439453125, 3951.03540039062, 
    3936.5751953125, 3936.5751953125, 3923.9765625, 4239.802734375, 
    4215.6904296875, 4293.3291015625, 4100.04736328125, 4293.56689453125, 
    4253.87744140625, 4189.19287109375, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 110, 472.108337402344, 
    1765.73474121094, 2963.14794921875, 3436.46337890625, 3443.97192382812, 
    3703.984375, 4150, 4150, 4150, 4150, 3721.27612304688, 2473.50634765625, 
    1478.68884277344, 882.745361328125, 1090.21459960938, 2009.16455078125, 
    3510.63745117188, 3704.70288085938, 3704.70288085938, 4150, 
    4385.37548828125, 4549.2919921875, 4719.65234375, 4642.2646484375, 
    4471.87646484375, 4552.51953125, 4605.1826171875, 4595.95458984375, 
    4432.83740234375, 4224.1279296875, 3998.60913085938, 3817.53515625, 
    3623.95361328125, 3395.4736328125, 3148.61767578125, 2800.80322265625, 
    3182.24536132812, 3461.03564453125, 3667.7626953125, 3897.57739257812, 
    3983.390625, 4034.06030273438, 4238.64111328125, 4369.990234375, 
    4403.50537109375, 4403.50537109375, 4641.12646484375, 4468.0927734375, 
    4391.90234375, 2538.25170898438, 2538.25170898438, 2363.06079101562, 
    3355.40087890625, 5012.63427734375, 5092.1669921875, 5153.50439453125, 
    5217.19189453125, 5034.65283203125, 4911.271484375, 4725.31689453125, 
    4299.81591796875, 3697.45751953125, 2998.1474609375, 1652.27990722656, 
    316.278015136719, 230, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 2559.19506835938, 2913.064453125, 2939.39111328125, 
    2702.75048828125, 2250, 2268.60327148438, 4969.8544921875, 
    4991.251953125, 4970.7060546875, 4859.17138671875, 4579.69140625, 
    3855.24194335938, 2018.6650390625, 2018.6650390625, 1937.41796875, 
    2157.224609375, 3065.78548661781, 4290.42431640625, 4720.81201171875, 
    4756.130859375, 4894.6767578125, 4891.26025390625, 4385.1884765625, 
    4192.001953125, 4390.302734375, 4390.302734375, 4220.5283203125, 
    4160.00927734375, 4125, 4235.95458984375, 4373.56298828125, 
    4550.283203125, 4675.75732421875, 4675.75732421875, 4562.419921875, 
    4532.84912109375, 4537.375, 4404.7353515625, 4385.6533203125, 
    4248.5087890625, 4240.8935546875, 3952.75708007812, 3822.166015625, 
    3318.89721679688, 2968.47338867188, 3163.19702148438, 3398.06616210938, 
    3405.24584960938, 3763.35546875,
  4000, 3908.30151367188, 4176.2978515625, 4213.1728515625, 3884.06591796875, 
    3726.12670898438, 3321.99337280395, 2067.52587890625, 2375.466796875, 
    2866.97192382812, 2866.97192382812, 3115.48413085938, 3115.48413085938, 
    2344.91235351562, 2635.71362304688, 2848.65551757812, 3166.84594726562, 
    3166.84594726562, 2191.85384798669, 3179.12182617188, 4176.94482421875, 
    4395.07666015625, 4507.98583984375, 4743.6962890625, 4874.34326171875, 
    4814.15234375, 5189.9951171875, 5147.90185546875, 5211.0595703125, 5500, 
    5500, 5470.67138671875, 4995.56689453125, 2393.78930664062, 70, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    90, 4579.8564453125, 4527.93896484375, 4296.8037109375, 3547.93823242188, 
    2450.390625, 2450.390625, 1678.93835449219, 1429.56237792969, 
    1229.91088867188, 1637.74096679688, 3021.62577171615, 3021.62577171615, 
    3021.62577171615, 1939.81616210938, 1528.16613769531, 2391.3359375, 
    2391.3359375, 2363.7021484375, 2690.83057001283, 2762.00390625, 
    3953.82543945312, 4261.74365234375, 4268.4775390625, 3980.58984375, 
    3224.76000976562, 2526.73046875, 2098.17529296875, 1935.05359591651, 
    3272.099609375, 5500, 5500, 5500, 4848.8408203125, 5500, 
    5436.84716796875, 5435.35595703125, 5467.39306640625, 5402.279296875, 
    5407.79052734375, 5458.13916015625, 5249.13037109375, 5223.41162109375, 
    5212.7392578125, 5317.927734375, 5275.41064453125, 5295.474609375, 
    5339.88232421875, 5081.80615234375, 4782.7158203125, 4923.2275390625, 
    4998.96337890625, 5020.93896484375, 5096.083984375, 5114.33251953125, 
    4901.00439453125, 4577.93212890625, 4341.0703125, 4676.8330078125, 
    4716.36572265625, 4707.92822265625, 4617.5546875, 4692.17138671875, 
    4659.81787109375, 4293.93603515625, 4167.4873046875, 4114.54541015625, 
    4180.38330078125, 4341.09521484375, 4119.4111328125, 4134.251953125, 
    4188.06591796875, 4234.77783203125, 4236.9384765625, 4204.998046875, 
    4158.06591796875, 4101.57177734375, 3978.2197265625, 3985.509765625, 
    4019.5751953125, 4007.87939453125, 3861.36962890625, 3745.89721679688, 
    3721.27612304688, 3705.30419921875, 3678.85546875, 3577.31616210938, 
    3503.52270507812, 3466.00830078125, 3414.44775390625, 3333.87036132812, 
    3305.39819335938, 3170.24755859375, 3046.67529296875, 2840.66748046875, 
    2875.9423828125, 2953.25756835938, 3026.07153320312, 3144.6513671875, 
    3089.2333984375, 3115.86083984375, 3115.86083984375, 3305.72509765625, 
    3439.93603515625, 3388.09912109375, 3439.83569335938, 3585.42822265625, 
    3369.59008789062, 3627.80151367188, 3633.60620117188, 3562.9991148724, 
    3690.3994140625, 3690.3994140625, 3606.19384765625, 3356.42529296875, 
    3345.23388671875, 3372.89526367188, 3501.21313476562, 3689.15991210938, 
    3885.40209960938, 3792.7568359375, 3755.89013671875, 3729.63330078125, 
    3865.69750976562, 3913.36596679688, 3942.97045898438, 4009.26684570312, 
    3876.9736328125, 3795.18115234375, 4201.52587890625, 4174.25927734375, 
    4025.90771484375, 4168.22265625, 4189.19287109375, 4189.19287109375, 0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 80, 130, 1221.5498046875, 2321.734375, 3387.2978515625, 
    3637.3544921875, 3703.984375, 4022.4267578125, 4150, 4150, 4150, 
    4261.60009765625, 4150, 3074.62768554688, 3074.62768554688, 
    2430.28247070312, 3365.7177734375, 3404.79223632812, 3696.28735351562, 
    3482.68798828125, 4150, 4077.42724609375, 4745.193359375, 
    4903.54931640625, 5130.755859375, 5045.9150390625, 4633.7705078125, 
    4494.79150390625, 4604.95458984375, 4472.8662109375, 4349.04736328125, 
    4111.56591796875, 3955.32373046875, 3826.35083007812, 3576.97290039062, 
    3529.4765625, 2927.81225585938, 3171.71850585938, 3576.30712890625, 
    3667.7626953125, 3979.29809570312, 3991.7734375, 4166.3447265625, 
    4125.67724609375, 4319.14111328125, 4403.50537109375, 4403.50537109375, 
    4660.72900390625, 4706.96630859375, 4482.28271484375, 4143.82080078125, 
    3695.72436523438, 2653.2548828125, 3389.2653479186, 5043.7568359375, 
    5040.6875, 5176.6103515625, 5234.9990234375, 4834.0732421875, 
    4941.4765625, 4703.98974609375, 4073.71240234375, 3578.33544921875, 
    2622.96850585938, 608.20849609375, 170, 170, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 80, 1565.60656738281, 2218.86865234375, 
    2429.91259765625, 1919.65515136719, 2358.80984022471, 4938.5556640625, 
    4964.916015625, 4899.771484375, 4841.439453125, 4679.083984375, 
    4190.5712890625, 3082.52856445312, 2450, 2453.50268554688, 
    2453.50268554688, 3154.52197265625, 3203.27294921875, 4209.9052734375, 
    4598.939453125, 5047.9716796875, 4903.61474609375, 4623.9482421875, 
    4707.955078125, 4606.71826171875, 4804.96630859375, 4902.83349609375, 
    4514.6083984375, 4159.38818359375, 4125, 4125, 4333.26025390625, 
    4435.35791015625, 4575.08447265625, 4557.8095703125, 4464.6572265625, 
    4419.18185522252, 4136.796875, 4140.5517578125, 4098.7001953125, 
    4130.06201171875, 3946.2880859375, 3410.09765625, 3294.46313476562, 
    3090.96142578125, 3434.97265625, 3590.21997070312, 4004.08056640625, 
    4000.32836914062,
  4130.04970597464, 4243.17088979408, 4218.25017509699, 4353.41919899949, 
    4194.91066908332, 4038.51037143336, 3321.99337280395, 2514.33457333003, 
    3065.78548661781, 4028.0642239222, 4121.27969268171, 4272.47111633591, 
    4138.07552418271, 3440.16294574566, 3148.18158392622, 3149.13801439716, 
    3988.84406886356, 3901.33223298542, 1465.08693161149, 3460.46023409179, 
    4265.62018975029, 4265.62018975029, 4248.60169220788, 4373.77544219693, 
    4753.62784698857, 4812.66458304871, 5228.34538225312, 5167.70344130337, 
    5360.74682660662, 5500, 5402.47375706515, 5287.89936811369, 
    2844.48899782977, 453.703763993212, 70, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 90, 2810.69578281359, 
    4200, 4200, 3547.93823242188, 2870.61777683132, 2870.61777683132, 
    2125.21936974611, 1595.91493594391, 1514.73977730206, 1539.02046072481, 
    3021.62577171615, 3021.62577171615, 3021.62577171615, 1376.65945425706, 
    2864.25522671102, 2864.25522671102, 2693.26209966418, 2693.26209966418, 
    2690.83057001283, 2910.18384813044, 3511.20993563703, 4014.21467715261, 
    4014.21467715261, 3899.71168206782, 3529.5283669988, 3269.07653100471, 
    1760.60122418777, 2056.49380264939, 1936.73584172348, 4169.73674027006, 
    5500, 5500, 3787.09595147351, 5357.47763546844, 5249.78073040947, 
    5031.45937341807, 5500, 5436.11617638433, 5191.08316505282, 
    5473.95459844324, 5500, 5199.0988177041, 5375.65871365297, 
    5133.1283413138, 5133.1283413138, 4732.87200157008, 5064.04349306078, 
    5041.10100797465, 5097.44847155076, 5072.05565367222, 5115.44483351133, 
    5085.14132368297, 5119.88133975654, 4891.88747125624, 4536.17630335457, 
    4613.24170319485, 4567.01067495847, 4746.82674353236, 4582.38137951942, 
    4337.04420605039, 4262.21543263798, 4222.38804800332, 3701.82089549313, 
    3426.50903037553, 3608.44194939128, 3608.44194939128, 3859.20567256003, 
    4271.0587602387, 4251.42201016258, 4157.72600032904, 4173.16348242766, 
    4162.36352644917, 4114.16151696418, 4180.98602672822, 4084.63701361757, 
    3882.70632799919, 3970.96777768374, 3985.509765625, 4032.38659972786, 
    3758.40335849289, 3722.53846736055, 3754.41932789085, 3674.04993790706, 
    3556.43885023192, 3531.27626718379, 3523.57188139583, 3343.88373848461, 
    3558.764375562, 3513.24118460263, 3278.84820118985, 3274.91797215046, 
    3079.03471696126, 3030.42376815261, 2852.52774025066, 2983.49139422074, 
    2923.85009396995, 2879.45810031449, 2989.98823566213, 3087.16024154015, 
    3077.38993453031, 3179.21667791772, 3305.72509765625, 3393.01002946419, 
    3423.94795518752, 3430.34847029756, 3510.91930793407, 3569.22038410294, 
    3586.19918947113, 3562.9991148724, 3646.87693402606, 3534.69975279694, 
    3699.87642012147, 3464.41146208422, 3398.74574283354, 3171.3616641935, 
    3246.57122143772, 3227.44518757928, 3439.00743878882, 3627.81777884548, 
    3654.84016429293, 3654.84016429293, 3788.89572341305, 3901.64174822343, 
    3845.03312898055, 3967.90846157093, 3942.97045898438, 3939.39416953128, 
    3972.28592751322, 3861.74403779221, 4025.90771484375, 4025.90771484375, 
    4202.35760188567, 4074.86111081024, 4074.86111081024, 1669.28501571787, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 110, 301.156558774663, 1979.4273033476, 2986.87187844271, 
    3565.59290618302, 3693.4508245992, 3286.52304345131, 4150, 4150, 4150, 
    4351.33855302784, 4214.63731726617, 4305.2024551374, 4295.11280295987, 
    4135.70792036822, 3651.79409179606, 3311.12484133135, 2888.92173901412, 
    3145.3054905966, 4150, 4719.56967597936, 4939.7932777188, 
    4996.70318885084, 4884.54444978891, 4919.07268000636, 4754.81421859496, 
    4674.15997819337, 4561.94542444473, 4507.49319292624, 4321.41414210246, 
    4302.41972251197, 4030.41078665484, 3913.84315494075, 3700.70159318108, 
    3411.97586830084, 3171.55170841943, 2868.80809725452, 3301.78449306327, 
    3633.36087507443, 3912.64164396276, 4073.15615224979, 4279.25794147504, 
    4340.18279274077, 4325.46236752036, 4453.98377684169, 4572.63993088596, 
    4623.69054246586, 4507.13454224791, 4551.76228018725, 4426.67669704125, 
    4329.64528757099, 3609.19561418435, 3389.2653479186, 4985.29602781583, 
    4973.47859606898, 5000.76434246508, 5037.0768100692, 4870.486043097, 
    4931.07800840881, 4703.98974609375, 4372.37468242229, 3688.51953272567, 
    2512.92784816316, 370.154968261719, 170, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 552.393538428005, 1820.40078752131, 
    1866.6905047022, 1919.65515136719, 2358.80984022471, 4529.76426063048, 
    4840.52988243793, 4780.95171281013, 4679.75126017681, 4568.61171330343, 
    4275.33409538548, 3916.52053744345, 2450, 2453.50268554688, 
    2453.50268554688, 2453.50268554688, 2438.30848177109, 4079.44832165225, 
    5077.62886582415, 5095.47338534044, 5126.46210686765, 5040.03104147857, 
    5021.60382945021, 4992.42033650029, 5091.71741473185, 5091.71741473185, 
    4637.56724002281, 4469.29631525392, 4176.80678156318, 4125, 
    3513.01180017582, 3513.01180017582, 3991.07425969921, 4332.1624062016, 
    4200.02295177138, 4271.46006596504, 4260.14230157586, 4126.65684669029, 
    3818.5343495561, 3799.41658926619, 3569.17291839313, 3387.2978515625, 
    3183.0885141089, 3392.67733428754, 3692.00626338207, 3675.69122551279, 
    3891.7847600419, 4000.15937717402,
  4065.89147763595, 4238.55967267988, 4229.54794514849, 4395.88128788579, 
    4367.50429404821, 4098.89904921892, 3543.87226324013, 2514.33457333003, 
    3469.00070806534, 4309.29080061053, 4691.20743626289, 4554.17075059391, 
    4298.68065454887, 4304.64381590663, 4291.46490016951, 4265.75546398614, 
    4371.49281251049, 4102.98362085469, 3467.59801067686, 4305.20418766379, 
    4547.05633411415, 4677.71132132096, 4629.1611353112, 4658.36793640569, 
    4799.89106125237, 4919.11363706249, 5262.6596735458, 5369.9392418888, 
    5305.05581976056, 5412.82695613091, 5143.41858983545, 3598.57938155268, 
    1290.26495406263, 425.785466617812, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 598.582848291803, 
    3688.85086219544, 4137.06277011802, 4137.06277011802, 3276.33298540559, 
    3102.61688041099, 2870.61777683132, 2177.03019929976, 1605.51794667436, 
    1492.88374562634, 1703.18479519602, 2952.8164921715, 3344.15361951335, 
    3217.40357434331, 1777.00088392329, 2864.25522671102, 2864.25522671102, 
    2905.69181851232, 2977.30818871205, 2891.96429881867, 3518.78967177782, 
    3899.24302456478, 4350.07296817072, 4194.05032445765, 4031.61764443499, 
    3794.67040679068, 3148.04258665972, 1731.15438875342, 2217.7497327348, 
    2259.04726938006, 3558.63092204947, 4272.28519789941, 4272.28519789941, 
    5151.13204937381, 5253.89301329408, 5143.41858983545, 5151.82807043689, 
    5484.59461161303, 5500, 5500, 5468.2582402431, 5500, 5449.8441988633, 
    5411.25574173621, 5342.96212595621, 5078.95139239648, 4984.48129841096, 
    5115.14285796601, 5023.87579437964, 5072.05565367222, 5072.05565367222, 
    5085.14132368297, 5085.14132368297, 5061.00903217242, 4835.7702891213, 
    4454.80516107727, 4095.33479009229, 4511.03202871705, 4461.92403644509, 
    4168.17952750381, 3695.52712363539, 3083.79958942393, 2244.17530361707, 
    2540.99217165055, 3387.2978515625, 3758.64637489801, 4014.96598682426, 
    4220.46866499158, 4326.91311333094, 4212.83271263619, 4217.32168431711, 
    4149.49769734364, 4122.52060134785, 4077.29020326625, 3993.0224086224, 
    3977.9313877401, 3955.65253503337, 3956.79231870643, 3899.67135514762, 
    3810.49705938271, 3808.16367928121, 3820.56925686961, 3688.45068004634, 
    3614.2904252827, 3491.17130815751, 3411.67607212435, 3347.90833360694, 
    3343.88373848461, 3374.03806710875, 3374.03806710875, 3266.80874890392, 
    3083.00401979317, 3028.00055473644, 2701.57027712264, 2665.09140644818, 
    2718.0926594849, 2718.0926594849, 2735.64383247666, 2959.34062931019, 
    2844.54085719189, 2836.18624917577, 2674.91589739519, 3018.66855827923, 
    3359.01792640043, 3270.38887406267, 3285.65821968378, 3222.63650452944, 
    3408.30452362822, 3442.44798329721, 3420.21470987184, 3396.7845816362, 
    3460.20711734538, 3545.65009136206, 3458.40625667329, 3612.21779441754, 
    3645.16301652947, 3686.02258906327, 3570.58160555255, 3427.26979091165, 
    3371.40702160615, 3683.27163665287, 3654.84016429293, 3823.68296182171, 
    3739.53673060724, 3846.04479196301, 3828.18094296334, 3989.87576763246, 
    3955.40969424004, 3822.06989672482, 4050, 4050, 4050, 4050, 4050, 4050, 
    3781.65701997948, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 347.285492451915, 1441.29322514436, 
    2295.31555450416, 2725.80635863034, 2851.45910506122, 2836.20427168033, 
    3172.29340131743, 4150, 4150, 4244.25490484775, 4265.69802044535, 
    4267.2096522141, 4267.2096522141, 4278.60099504976, 4356.87893571387, 
    4431.62046959384, 4566.90825442193, 4735.15880382443, 4820.43450339191, 
    4905.99706206238, 4964.2896881696, 5010.90815830123, 4883.19860953033, 
    4874.6928348152, 4837.27410790798, 4700.81410964451, 4659.6063970409, 
    4447.25196763893, 4368.06375002399, 4188.79402077313, 4025.36923166822, 
    3792.07810227472, 3583.97934276751, 3404.69051131505, 3111.3684889767, 
    3344.24163557876, 3438.97347823814, 3648.15779103425, 3898.32448331561, 
    4146.71276469288, 4139.97651769806, 4345.64720085662, 4360.12540549873, 
    4467.34565836146, 4627.41712027848, 4673.3199122047, 4688.22175845735, 
    4756.17854801362, 4720.784670925, 4561.77610212979, 4162.34550615586, 
    3193.54849468975, 4240.82988252286, 4524.56517260274, 4782.14816378248, 
    4870.486043097, 4889.32581648231, 4850.912164561, 4659.54947549622, 
    4357.45823504103, 3556.20361620099, 2101.23232371475, 713.645284248567, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    1354.54550139175, 1548.75423199767, 1737.94963000608, 2191.85384798669, 
    4194.13998706414, 4510.86430305793, 4615.896971949, 4551.3969743444, 
    4422.31085390515, 4275.33409538548, 3908.16321250272, 2230.97292955744, 
    1963.44369222536, 1678.01086309505, 2381.39282189074, 3249.90067386452, 
    4661.57728085578, 5115.1290585818, 5287.53687622229, 5299.65856060897, 
    5301.49005651965, 5143.41858983545, 5094.60213311098, 5102.90223778457, 
    5223.45183734046, 5255.26570808033, 5115.05526891491, 4864.39442626429, 
    4427.15875153804, 4137.18005886292, 3791.78318194838, 3721.27612304688, 
    3829.12661866819, 4000.85835133454, 3750.76416004187, 3897.81694861604, 
    3808.30523154608, 3637.14945091668, 3433.29189913431, 3209.82770902734, 
    3194.89645320192, 3321.59767393036, 3600.41446066078, 3817.65929639173, 
    3779.91925488157, 4038.84296649908, 4035,
  4170.63108524582, 4221.25016457579, 4324.57551060707, 4373.43953297949, 
    4373.43953297949, 4160.31669458408, 3453.25444216436, 2514.33457333003, 
    3622.78802782165, 4407.20919616552, 4794.73987800048, 4783.61568260597, 
    4606.59494575004, 4582.30535610321, 4578.8788839918, 4644.03912636511, 
    4747.72913184857, 4747.72913184857, 4677.4490478961, 4268.69275965733, 
    4451.97651712323, 4695.77498149507, 4928.33072104389, 4935.35679696171, 
    4902.17092342198, 4977.66879562253, 5047.37142701511, 5047.37142701511, 
    5125.79345030561, 4648.15942530949, 3855.13603187726, 2232.00546399652, 
    1033.56580065904, 70, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 1200.62896893604, 3688.85086219544, 
    4216.41764683475, 4236.84470010854, 3292.03305172377, 3228.21828543352, 
    2341.30588940991, 1923.0417239584, 1567.72921817894, 1512.5939183985, 
    1835.94180849488, 2732.19145868561, 3184.71274960557, 3085.52802787989, 
    1939.64875781125, 2546.44385381085, 2797.63493384722, 3009.53947639045, 
    3558.32932359464, 3707.10698831117, 4021.89530155629, 4231.13330321053, 
    4405.66231415225, 4324.9340008769, 4140.66316947843, 3813.15483243059, 
    2857.01927011859, 2221.61015767072, 2217.7497327348, 2238.54970057615, 
    3073.19527751297, 4342.66175275086, 4403.50400951895, 5235.57864459612, 
    5290.27175486947, 5374.50155693674, 5461.96325184829, 5499.9236655526, 
    5500, 5500, 5500, 5485.02746400498, 5419.4819106827, 5424.15827777244, 
    5332.43998569524, 5078.95139239648, 5024.0560859724, 4993.950563962, 
    5028.67390019976, 5098.49902274328, 5081.70617500708, 5056.40638745122, 
    4930.24490946628, 4815.59862110962, 4744.78114736523, 4589.27742967214, 
    4310.5735256199, 4310.5735256199, 4255.4920916757, 4011.47728558016, 
    3099.95499474951, 3316.42245533443, 3568.87113275539, 3801.30120072225, 
    3835.34257729635, 4097.02750933481, 4270.06951907413, 4279.73748110154, 
    4238.90201279945, 4228.37149208108, 4210.04531963034, 4190.88081634226, 
    4134.22810628455, 4014.88330681784, 4008.84541463564, 3856.96419652146, 
    3728.15245708428, 3721.27612304688, 3780.84486000863, 3755.4331640747, 
    3724.76118387482, 3679.32319007998, 3643.76654085545, 3548.14482693473, 
    3406.15604975124, 3333.7267574288, 3291.18080643427, 3271.9346200235, 
    3231.75708311619, 3151.7371098196, 2927.68259070678, 2878.09162672127, 
    2784.59103884648, 2885.86153966193, 2782.76144572558, 2849.21872312184, 
    2934.38388572984, 3104.53882587139, 3112.3747571286, 3040.20332568657, 
    2758.41088867188, 2723.48749954695, 3070.49278240527, 3065.78548661781, 
    3067.98102796027, 3142.34158947543, 3051.18084700638, 3327.43907723542, 
    3436.82809905361, 3446.53583689279, 3332.12940522169, 3282.60789787486, 
    3444.34263788113, 3389.6458777007, 3268.9583629368, 3560.36507022261, 
    3499.56953493758, 3491.8637225317, 3480.66220545118, 3358.92701208747, 
    3356.73577467507, 3544.322006658, 3698.74487833286, 3704.52075558775, 
    3704.52075558775, 3742.30619430216, 3902.54273761764, 3780.35033539675, 
    3892.25272968249, 4050, 4050, 4050, 4050, 4017.65260950183, 
    4039.09998658205, 4039.09998658205, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 334.244736680591, 
    673.168189330021, 1555.76596340374, 2172.35627711298, 2368.49020948947, 
    2534.54644236146, 2745.82558520821, 3228.30730916764, 4027.59887178456, 
    4027.59887178456, 4265.69802044535, 4353.89686204892, 4395.94625696463, 
    4443.47178735976, 4452.12593823663, 4561.73325522178, 4884.3308481158, 
    4983.33264264742, 5098.20034132639, 5083.13536366454, 5120.60625640023, 
    5025.3054174596, 4992.81193645737, 4869.6209307359, 4800.20269873261, 
    4647.20733351532, 4637.75511377971, 4448.82816998867, 4357.05107396864, 
    4175.40028432296, 4084.52017050723, 3868.11347537232, 3584.64129337209, 
    3339.99222163381, 3187.71400875199, 3431.17212859253, 3676.31652514003, 
    3887.97048883937, 4055.35771753258, 4088.65023279901, 4247.65964020839, 
    4402.51483664531, 4469.09720707317, 4576.13714781562, 4666.66629670527, 
    4768.57438033915, 4843.83792636489, 4949.06391161969, 4920.23541517288, 
    4709.89596466775, 4523.05543945419, 3638.86107614402, 3262.30444769182, 
    3082.59495940385, 3901.37923204169, 4595.5971585084, 4733.15526618951, 
    4744.26430848736, 4483.67088367407, 3987.29624818454, 3036.45985630902, 
    1548.13285289387, 707.791336663412, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 860.34900699956, 1170.90527014303, 
    1671.32455582663, 2310.35585059744, 3721.27612304688, 4189.28859554725, 
    4319.15775808308, 4349.48370510366, 4251.6030949895, 4003.5939036041, 
    3430.98177416991, 2230.97292955744, 1768.1383575229, 1678.01086309505, 
    2834.25610112025, 4006.6760744058, 4677.21208992919, 5059.9947969076, 
    5198.58510168983, 5270.33821557672, 5242.03840444192, 5184.3618920597, 
    5123.63718856849, 5102.90223778457, 5210.24892546068, 5189.25905013667, 
    5115.05526891491, 5088.00524958576, 4785.43652682823, 4516.82085763071, 
    4400.24103372465, 4228.04405739572, 4184.04022336469, 3897.58821250629, 
    3749.8918757941, 3579.31464526711, 3518.00908059251, 3377.20526304306, 
    3242.57927199852, 3199.7467826794, 3329.18592699495, 3581.7165112426, 
    3721.27612304688, 3936.64936076732, 4001.56517226959, 4047.48611341481, 
    4038.84296649908,
  4129.62025594702, 4245.06544615096, 4342.57118820929, 4377.74385711509, 
    4385.63366066429, 4192.74722935635, 3758.92241697352, 2450, 
    3688.54054756258, 4468.7286119359, 4787.55185638068, 4846.11832208212, 
    4810.13311482503, 4842.96027710625, 4892.42549406734, 4979.91781596674, 
    5079.96969847571, 5097.50415185396, 5069.0660909329, 4758.28218878442, 
    4093.58856317153, 4658.90457869435, 4964.90795224914, 5059.1757519723, 
    5042.62265314627, 4946.07482992966, 4810.51924430932, 4705.52119903163, 
    4382.53736220073, 3919.63486202158, 3205.77769859713, 1938.62990581942, 
    958.639324409817, 70, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 1517.27347491937, 3439.74884767343, 
    3813.60956119365, 3866.1835018099, 3292.03305172377, 2846.10213327557, 
    1992.18009779946, 1836.5015293951, 1545.26875627066, 1577.50262982867, 
    2074.08422846403, 2704.20555730691, 2790.83174201673, 2790.83174201673, 
    2140.62836982014, 2259.40807657782, 2572.00310639395, 3009.53947639045, 
    3698.94733047918, 3971.22193744431, 4205.89183421572, 4380.47619149948, 
    4333.42854817502, 4376.93669443876, 4159.89232599685, 3674.46409453601, 
    2772.53255115215, 2233.09358475916, 2083.89254584475, 2097.73825211526, 
    2498.38487354641, 4342.66175275086, 4982.24403052868, 5329.39034316341, 
    5441.55013960065, 5500, 5500, 5500, 5500, 5500, 5500, 5489.54122977282, 
    5428.83788679287, 5366.93523121161, 5249.28100822058, 5032.4212490823, 
    4986.59976560915, 4973.57611019054, 4961.20766762177, 4950.37987965817, 
    4908.53131928046, 4895.0179319176, 4795.05158749994, 4686.68112643318, 
    4610.79516303237, 4506.86440078033, 4310.5735256199, 4310.5735256199, 
    4312.32491330413, 3994.39450597886, 3660.74820050267, 3780.26054763866, 
    4036.1731480386, 4176.56842232826, 4252.22572767252, 4306.90184311616, 
    4336.73203499361, 4307.23682568614, 4193.086257612, 4205.18076833969, 
    4162.74251119982, 4102.3493201746, 4009.957024093, 3967.12604520287, 
    3905.76829935057, 3787.17191112393, 3694.36846799669, 3564.45119646804, 
    3583.84977303869, 3538.59699312402, 3522.07405543561, 3475.51365592755, 
    3425.41517804518, 3387.30621995946, 3299.27101266061, 3194.48104256381, 
    3079.12518772046, 3097.74659857904, 3085.5618224434, 2905.40155920799, 
    2898.75829614332, 2979.07961496354, 3018.98675171447, 3037.10745337034, 
    2973.11183944416, 3028.99978528837, 3185.62925272638, 3305.71204962413, 
    3376.67253247949, 3322.35718737023, 3375.15916425367, 3346.20858814425, 
    3260.19356291725, 3282.85383530423, 3327.28419679483, 3183.5637369676, 
    3170.25449985619, 3040.22998237743, 3274.28939017299, 3262.09116135402, 
    3218.47964423569, 3306.56564742617, 3285.82432745714, 3220.32218758882, 
    3212.46920573561, 3299.96884761102, 3328.82237874485, 3328.82237874485, 
    3328.82237874485, 3319.27714081661, 3340.37059109061, 3070.25116963963, 
    3339.05425814481, 3351.2507939702, 3351.2507939702, 3756.43300589855, 
    3952.41630438794, 4111.88086887032, 4088.40194803055, 4050, 4050, 
    3749.78539601327, 3948.38134735866, 4039.09998658205, 4039.09998658205, 
    4039.09998658205, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 240.561416625977, 460.795415826947, 
    751.84451263033, 1531.37201060798, 1893.14334134199, 2138.52732260812, 
    2527.33609525053, 2988.49735159664, 3491.97950407711, 3898.61157036895, 
    4097.23423570347, 4229.62601326259, 4289.0997683235, 4488.96259580082, 
    4651.52180065304, 4806.46262937177, 5037.30745591176, 5188.03072086498, 
    5240.94112322561, 5259.97898137901, 5229.84744278434, 5129.05905861854, 
    5045.71489070029, 4930.74193997593, 4828.41365506694, 4684.97556167094, 
    4597.66494915089, 4526.19373947857, 4356.81594105931, 4186.09024995742, 
    4106.78513248386, 3922.51643824655, 3695.19666110263, 3407.81504016227, 
    3344.11973632775, 3483.28858533049, 3708.08379061909, 3965.47203723904, 
    4175.40501265917, 4380.14547090418, 4460.916018357, 4568.94654364787, 
    4659.35978094293, 4761.36297775296, 4840.76382569532, 4942.54071364061, 
    5008.62360957119, 4997.67061054745, 5075.54137272006, 4992.18084313171, 
    4726.61029810396, 4390.48450794376, 3830.30230814673, 2970.66908088546, 
    3076.03688086331, 4041.47395704149, 4493.72147358842, 4534.81508565769, 
    4286.55722169857, 3684.04164187872, 2758.41088867188, 1478.68884277344, 
    730.099028488691, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 580.953491210938, 813.783205142792, 1485.19614601662, 
    2261.83768809263, 3120.64406627867, 3617.24588998514, 3903.67290891671, 
    4029.50018006597, 3969.97483317296, 3751.96959459619, 3252.46912358287, 
    1697.12502302956, -0, 1539.52340788021, 2916.26316166098, 
    4006.6760744058, 4543.03905844656, 4936.61665334032, 5085.91521683377, 
    5098.89821975592, 5066.16325136943, 5021.83824839001, 4974.6770050089, 
    5032.10030354546, 5084.06164940445, 5108.12056144014, 5062.08514591651, 
    4925.57469274506, 4811.59885021003, 4645.73039003495, 4400.24103372465, 
    4307.53805682028, 4142.85030612649, 4022.75619891772, 3807.12224909431, 
    3539.14141350261, 3341.45923198451, 3236.29861421444, 3327.21939115067, 
    3429.22920404735, 3529.01099674852, 3780.98126382114, 3900.20090723003, 
    4043.47382623819, 4101.36345772905, 4208.73033156926, 4143.63704676482,
  4275.98935025516, 4319.91165998098, 4366.61699642038, 4377.74385711509, 
    4377.74385711509, 4215.63011855828, 3900.40906239898, 2650, 
    3934.64679458308, 4528.14010036148, 4835.59118942226, 4935.99101762941, 
    4909.22623960055, 5021.23730650222, 5074.77224408145, 5143.84350440161, 
    5241.3124377265, 5309.10684695882, 5314.19616327954, 5218.95397584822, 
    5035.14544062991, 4855.22146940084, 5014.59802563496, 5066.59214559651, 
    5017.64120857399, 4837.5342151758, 4710.70331998565, 4068.52991343902, 
    3741.88212276044, 3683.95051507361, 3151.81238207084, 2074.06537861684, 
    1238.34590443145, 70, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 658.602779396555, 1517.27347491937, 
    2903.64551362136, 3028.81260543643, 3028.81260543643, 2801.92744448877, 
    2532.71888671197, 2051.35268642626, 1778.98973086404, 1592.31104336679, 
    1712.72500893013, 2281.8964709166, 2709.54742473887, 2704.20555730691, 
    2528.93906782579, 1990.65811859568, 2158.0596135651, 2536.79454952133, 
    3247.09169921523, 3710.85764481148, 4035.48888497929, 4194.01840454916, 
    4333.42854817502, 4396.0962821422, 4331.03627323711, 4094.64625024203, 
    3636.64523974662, 2852.88774966492, 2214.1180047755, 1882.37550796932, 
    2116.85258371872, 2559.77458095327, 4287.43964770477, 5143.41858983545, 
    5499.14550445891, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5456.29968890867, 5251.49930511239, 5253.98393836866, 5101.44873503467, 
    4977.26986497824, 4900.32426637085, 4847.54385597227, 4811.23770013371, 
    4826.44806402904, 4763.68574482341, 4758.0495103006, 4703.71668982256, 
    4666.55564144917, 4581.33595354001, 4525.42956675091, 4541.18480584962, 
    4310.5735256199, 4121.90219910085, 4098.35934255726, 3989.05584234131, 
    4116.38944555794, 4300.19262167919, 4419.18185522252, 4454.59753289808, 
    4461.70777357378, 4381.79717364862, 4320.86518894141, 4198.81820139652, 
    4161.20432817571, 4065.89147763595, 3986.72137130287, 3898.87425152437, 
    3852.19966627968, 3777.11147445946, 3644.70881009564, 3559.41478727432, 
    3501.78658209209, 3394.36283372164, 3454.43574880596, 3398.08956585473, 
    3376.20127971063, 3248.58942354451, 3283.02182576871, 3300.06445473908, 
    3266.24128787454, 3232.15441111159, 3208.49607855068, 3157.67421994142, 
    3038.63444521911, 2985.35405876951, 3031.75073363399, 3132.67279892876, 
    3194.67596938187, 3178.8524707237, 3191.6926957011, 3366.04445839408, 
    3493.0244445173, 3564.1513864241, 3603.17882820958, 3582.14862570139, 
    3560.38831824842, 3559.5476906943, 3547.55764387319, 3520.9494228923, 
    3474.37276080145, 3453.86280772631, 3394.4447770916, 3449.50519132316, 
    3478.27671952432, 3497.13167652549, 3528.90310450301, 3454.43010819289, 
    3533.94499896027, 3576.23899668114, 3619.93511973014, 3556.50591917423, 
    3632.49712635151, 3579.12739340648, 3529.56232000675, 3596.32636570643, 
    3416.71245352087, 3441.09936969761, 3460.76394046813, 3540.83643613515, 
    3818.48993036311, 4048.41771647607, 4218.70556674742, 4300.38885025196, 
    4288.46468836507, 4215.86432920475, 4122.64809252176, 3887.95325757591, 
    4083.38731899196, 4172.20302241556, 4137.4537521979, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 299.674571381543, 506.525611873329, 831.355340372086, 
    1281.8531028924, 1697.12502302956, 2123.86310271776, 2647.85260545679, 
    3175.78926161887, 3634.97037425038, 3942.29725107297, 4126.02433065169, 
    4265.7784588929, 4462.11519806451, 4657.38738343252, 4871.47570811512, 
    5082.56453247434, 5210.34693318396, 5299.73658698268, 5351.40951058892, 
    5339.75276603559, 5305.44627513318, 5180.23748790566, 5072.68657754738, 
    4957.40785336838, 4865.20291463239, 4745.24695653404, 4583.22797882715, 
    4438.04248260875, 4324.88327771788, 4196.89241865499, 4011.18262920893, 
    3779.94673687141, 3550.16882392397, 3364.94763611858, 3463.21757726273, 
    3708.08379061909, 3968.06081556186, 4228.16014389579, 4425.1871074728, 
    4583.60802507453, 4678.73638680486, 4787.48344196823, 4884.36230117052, 
    4980.46544925369, 5031.24227423723, 5095.74349971937, 5132.79942088851, 
    5132.79942088851, 5114.82256871465, 4901.64197549331, 4493.64969544535, 
    3776.54812285271, 3027.00366799113, 3000.47014071994, 3762.35916667622, 
    4255.79054021911, 4351.11297703982, 4000.00917536216, 3335.85168545681, 
    2420.94524484664, 1341.82002836157, 685.151404079313, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    1326.24635387602, 2237.86162866415, 2919.43353882474, 3288.75733625709, 
    3532.00846194744, 3611.57563753279, 3593.44607799006, 3411.80210074478, 
    2855.52774441814, -0, -0, -0, 2466.66776221529, 3786.84460104126, 
    4342.20611259389, 4761.62668362541, 4932.57916636208, 4962.7678588968, 
    4865.78041171435, 4787.52335666941, 4794.83215699253, 4838.67529131632, 
    4907.21522880616, 4916.98873089652, 4858.07127730467, 4759.80855415892, 
    4611.29406054407, 4499.09345309135, 4387.98190728403, 4275.70742576829, 
    4084.34535140581, 3914.4348823189, 3670.32178770878, 3466.37760074827, 
    3257.58638447822, 3290.64871459137, 3405.85758805152, 3555.95267068187, 
    3721.27612304688, 3863.02562139269, 3996.63832349954, 4099.25139122234, 
    4167.44652450554, 4220.30487513238, 4277.63414055145,
  4406.93909432159, 4435.02686853828, 4451.45386865219, 4474.28237353917, 
    4447.89170885671, 4247.90518209934, 3962.91059225322, 3333, 
    4150.18552315763, 4572.80739470807, 4873.43084610599, 4967.7941700266, 
    5017.73018106873, 5089.03854170738, 5146.58431220602, 5205.90911594463, 
    5328.36144466083, 5449.42361945718, 5488.36130286214, 5405.03415320444, 
    5287.88132948114, 5061.59915796591, 5003.0010067476, 4954.42487622574, 
    4795.93916438524, 4727.37058303913, 4505, 4034.88084437255, 
    3740.06849018172, 3771.87116266214, 3592.9860366021, 2871.9832094614, 
    1829.70715672165, 1088.68810450859, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 190, 658.602779396555, 
    1295.84009271083, 2550, 2550, 2550, 2411.9314192889, 2249.00670817428, 
    1988.65620342361, 1813.12568372434, 1648.3371664196, 1956.54665472741, 
    2377.77027707637, 2665.34001729425, 2729.78766551144, 2266.29221078739, 
    1860.8553952277, 2113.31433636761, 2482.77334293811, 3247.03841881874, 
    3710.85764481148, 3967.04612358226, 4038.66114905438, 4121.35523906247, 
    4191.0451842763, 4187.23107890345, 4024.32240626634, 3591.67535905953, 
    2917.29114032725, 2295.53476379113, 1935.05359591651, 2164.21662224033, 
    2569.30806074812, 3884.62436079194, 5179.73235014496, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5407.89515994579, 5232.8009329998, 
    5143.81672107376, 4974.40061415652, 4849.41200315916, 4759.05532761955, 
    4711.07171051427, 4721.31721448639, 4744.56647367292, 4731.55935401327, 
    4709.80831856274, 4613.53066128589, 4553.2805203336, 4524.71990522333, 
    4487.44717502968, 4419.18185522252, 4279.8568570872, 4369.88811917926, 
    4197.80275837181, 4283.78385999065, 4363.24596905814, 4464.61598832407, 
    4539.56182337733, 4529.05211216299, 4472.27495879848, 4342.67734936369, 
    4235.26340090534, 4129.9435375496, 3960.68102447184, 3870.62770016362, 
    3761.88843965289, 3685.48249506229, 3707.83768875721, 3629.8478443261, 
    3534.00411914892, 3468.54722009487, 3479.82760177972, 3494.37923291359, 
    3535.94852651972, 3513.62374122156, 3499.54049174449, 3462.71025029994, 
    3434.98681085331, 3396.45116402431, 3362.90057838965, 3324.79821495051, 
    3307.14538134871, 3256.15479247201, 3175.27785631278, 3110.72844127508, 
    3096.53091268744, 3177.875706514, 3274.25682525982, 3316.96329564987, 
    3345.04434725698, 3480.18537777292, 3585.56902449894, 3682.442084854, 
    3729.51891510576, 3753.03971326393, 3755.51867336499, 3757.92194457467, 
    3753.26425970322, 3741.89966980278, 3705.90089559694, 3705.90089559694, 
    3694.35276721458, 3721.27612304688, 3728.14368728537, 3731.36445287934, 
    3703.90413972107, 3696.16936722349, 3709.12784613846, 3755.19335761301, 
    3822.53061894471, 3862.03982443479, 3884.94426426172, 3870.80491164601, 
    3798.84060931009, 3737.37406659968, 3594.10734053, 3517.43031518652, 
    3470.29686349246, 3529.67898846244, 3782.49098914998, 4033.33319084532, 
    4323.23279783555, 4461.95544191158, 4472.25512601052, 4376.07170450348, 
    4295.82359325192, 4128.50347785241, 4135.0542704557, 4137.4537521979, 
    4137.4537521979, 3146.80193254396, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    528.424953645431, 730.332413158285, 1043.12608339423, 1462.21416126929, 
    2238.62572908916, 2837.44639239522, 3352.11513329302, 3783.16642355822, 
    4065.89147763595, 4233.91482694526, 4399.28161801747, 4602.00867315233, 
    4824.20795668429, 5008.45638601948, 5177.11909808497, 5298.68327503892, 
    5373.70544323758, 5400.65110680117, 5374.24774888817, 5314.433325256, 
    5219.09869317235, 5121.22368388109, 5005.18336912404, 4846.7337372745, 
    4687.5760916545, 4567.6676325881, 4444.31542415121, 4307.04045454281, 
    4103.32646811808, 3863.16608458619, 3631.56691127524, 3461.81909341827, 
    3502.02150164264, 3705.5293506168, 3949.35266504641, 4244.03413133263, 
    4421.19842195965, 4580.10513059933, 4740.79253875101, 4875.57813015251, 
    4948.6799092277, 5038.15820345906, 5127.10861505736, 5176.39557014426, 
    5237.58312041057, 5244.10572975435, 5185.55939654447, 4982.88943208861, 
    4523.6487142817, 3766.67447002004, 3166.26203275163, 3148.41674795964, 
    3700.92151134836, 4016.95078107402, 4016.95078107402, 3756.56661793474, 
    2972.98458542247, 2070.62997047906, 1164.80634003826, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 570, 
    2179.16191045429, 2731.49615807304, 3065.78548661781, 3288.81309470592, 
    3325.05003294338, 3293.02991778292, 3093.91105496691, 2511.10764448436, 
    -0, -0, -0, -0, 3488.64426753851, 4079.48727263566, 4524.14568632179, 
    4796.79974581409, 4805.68201245752, 4670.88274523131, 4498.14491272971, 
    4467.46050804411, 4582.3856378491, 4669.28673375228, 4714.47645801227, 
    4634.14182325243, 4542.13646069301, 4419.18185522252, 4324.53339621404, 
    4213.37844295523, 4088.1584131897, 3952.96503519651, 3790.60141895392, 
    3560.76254526607, 3344.47182330956, 3232.06492824651, 3364.35090344665, 
    3533.67129541239, 3743.63233878803, 3879.81457844077, 3984.6379076075, 
    4094.841915681, 4194.76946688048, 4304.66623524972, 4336.52415989829, 
    4389.29479046407,
  4586.16912326963, 4585.57592051546, 4596.33844518516, 4579.03785739764, 
    4516.9549034989, 4304.27632703959, 4038.13130339401, 3333, 
    4174.44304876521, 4573.55438152792, 4845.03743391474, 4945.10307816789, 
    5019.43919363506, 5102.01078795585, 5168.81639224842, 5213.88948659803, 
    5346.74867597832, 5500, 5500, 5500, 5500, 5241.32396563711, 
    5048.91417399402, 4801.16730677605, 4505.02153913166, 4508.1009686592, 
    4505, 4126.07069597084, 4116.65072752822, 4156.2191538562, 
    3973.44590025259, 3451.46692046743, 2442.39054054829, 1478.68884277344, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 190, 555.872542718758, 1042.65290128262, 1710.68891456632, 2550, 
    2550, 2129.73637144263, 1996.03949780786, 1797.32250068938, 
    1764.26824652923, 1777.11606508842, 2057.68832792079, 2353.4608831765, 
    2639.5843222398, 2487.30482030053, 1953.63620684299, 1867.08925629296, 
    2134.30644933817, 2665.24685306533, 3283.84592561678, 3396.29238888299, 
    3554.89183421369, 3670.38345235014, 3756.07420334438, 3865.10367045026, 
    3917.65623736052, 3845.16919286788, 3535.08947987053, 3009.00004088572, 
    2390.30980293918, 1987.41070769959, 2150.90887168795, 2494.5729255217, 
    3261.2030859254, 4781.90185538265, 5430.74431834156, 5500, 5500, 5500, 
    5500, 5500, 5500, 5474.41317282213, 5346.23127504002, 5196.25894496046, 
    5044.98398327715, 4878.93115185147, 4763.1835070218, 4669.91888034256, 
    4651.50064518762, 4646.16037413862, 4671.45525074954, 4688.59021142698, 
    4647.44577165254, 4583.68364186514, 4497.9797336883, 4435.35137692775, 
    4328.91259463312, 4405.40111360637, 4430.92942303256, 4460.77599226567, 
    4466.08797615055, 4468.48970541947, 4446.04620269448, 4443.51423610024, 
    4478.84595944019, 4442.97081517397, 4368.65388678934, 4233.20227411648, 
    4041.54102303604, 3864.72238026479, 3776.70029276475, 3707.05428916106, 
    3639.21510044772, 3561.41798926813, 3569.88568235328, 3564.61592417846, 
    3549.73257437854, 3555.5973752015, 3595.49819880031, 3660.21941415773, 
    3706.08349818874, 3691.27638470446, 3661.03295728959, 3611.88199392496, 
    3554.20726141789, 3500.40407661416, 3443.41988952482, 3420.14170457373, 
    3395.4934602466, 3346.12348862643, 3266.93762069733, 3204.20731755884, 
    3191.18033694748, 3206.76911260621, 3281.46485354402, 3353.61624568471, 
    3445.22710520542, 3539.95102537927, 3639.49038328409, 3729.92945303298, 
    3794.0188376894, 3827.30234633426, 3846.98783421398, 3865.4087615103, 
    3885.05616879989, 3903.46544526408, 3902.63260084172, 3913.38048889897, 
    3901.45051146128, 3899.39169848062, 3892.88178931142, 3907.68156997911, 
    3898.45620076481, 3879.36514922968, 3886.71077782078, 3919.47503317499, 
    3984.25015710583, 4042.67518634029, 4047.12411285674, 4037.30824028639, 
    4006.2538864601, 3966.40749437145, 3880.08758524602, 3743.98449185722, 
    3501.15583828067, 3387.2978515625, 3599.70830882247, 3951.42039106625, 
    4312.37774179524, 4525.37390514703, 4592.10454533704, 4545.31782940758, 
    4469.33566133105, 4344.41682849833, 4319.78839039081, 4148.97844648417, 
    4379.52450888098, 3465.02072196186, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 1085.05843356077, 1697.12502302956, 2452.13869943843, 
    3025.62160107718, 3507.92626627224, 3886.79350424502, 4123.50655248632, 
    4313.32719334855, 4483.73628149263, 4661.52801887447, 4850.69265527823, 
    5046.00872212362, 5211.54361750208, 5309.31643440427, 5391.302169467, 
    5399.76517496048, 5353.02505031957, 5278.09512555725, 5185.39869434248, 
    5099.75676842587, 4965.819047089, 4826.80174110346, 4689.41767868348, 
    4544.6624840565, 4367.74225941342, 4167.31795217251, 3990.52203781764, 
    3765.31725041649, 3567.85546219026, 3512.69454141378, 3622.24239473013, 
    3859.62395981216, 4123.91299924795, 4353.87709188741, 4581.40192111753, 
    4748.21242290072, 4859.35636176266, 4961.88295165354, 5061.03229609622, 
    5143.41858983545, 5189.73316980975, 5254.93106950075, 5316.81449419577, 
    5253.92989331445, 5053.75552338893, 4684.94478453477, 4073.93021811718, 
    3483.65372826982, 3290.08412833393, 3537.22039957519, 3811.83929038399, 
    3814.40537176407, 3387.2978515625, 2635.73188916564, 1792.67801968854, 
    1016.28561289622, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 1199.58146437838, 2049.81531575107, 
    2622.05117528737, 2945.27758316167, 3095.46131385416, 3078.14718123661, 
    2994.42389570561, 2760.01279092483, -0, -0, -0, -0, -0, 3251.21094112802, 
    3966.66579155766, 4427.84896594736, 4713.63705314985, 4692.66749527368, 
    4495.7722330907, 4315.27649955633, 4237.33518508171, 4302.32540948322, 
    4408.81080887101, 4458.14414866975, 4428.99199356759, 4343.75121032504, 
    4221.93818718823, 4097.74422226575, 3978.09992097544, 3874.66480849105, 
    3745.83172987669, 3568.35043548301, 3361.65507262617, 3201.70257579734, 
    3193.40915115792, 3367.6332484637, 3631.96807252137, 3873.3160155477, 
    4016.39851864994, 4102.51730123787, 4207.95706380502, 4273.44958906613, 
    4387.82675381612, 4483.17088394398, 4552.63937651413,
  4736.77472323068, 4736.57767650498, 4740.51056791939, 4703.2639020272, 
    4589.45185795149, 4331.53195868943, 4024.89491363747, 3333, 
    4065.89147763595, 4486.55223748062, 4768.7159496115, 4919.37900985824, 
    4994.53678216462, 5070.29498002577, 5160.1002944529, 5218.67972425055, 
    5360.8784220364, 5500, 5500, 5500, 5500, 5449.57633004648, 
    5128.85585583997, 4663.87121450909, 4431.11385217117, 4575.96759786076, 
    4589.27977596717, 4419.18185522252, 4438.043721817, 4430.98220858166, 
    4149.18913610704, 3540.9055834814, 2442.39054054829, 1548.11043215947, 
    803.625015916513, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 110, 230, 545.419436106388, 1051.69511197961, 
    1803.19972842396, 2550, 2550, 1890.82155709655, 1774.92296151271, 
    1649.49011671483, 1753.05817372212, 1846.68562116194, 2044.67879189348, 
    2353.4608831765, 2353.4608831765, 2290.50571318798, -0, 2111.20707693595, 
    2336.38410883367, 2695.50666974581, 2963.61371914122, 3088.78793573769, 
    3209.9032991091, 3174.46949957337, 3231.95229602848, 3352.69145893815, 
    3545.47350335499, 3634.25933915523, 3445.96962237104, 3016.14950357872, 
    2414.73345596945, 2030.89247188587, 2033.64910367341, 2293.41136542742, 
    2816.84885311515, 4065.89147763595, 5233.76020129616, 5500, 5500, 5500, 
    5500, 5485.9217461387, 5452.12407729264, 5388.31223009016, 
    5276.65247915195, 5149.29628623736, 4999.58220832841, 4852.87868175799, 
    4729.24166645864, 4635.09839641065, 4554.21542494894, 4558.09434332041, 
    4575.41165153652, 4618.20603630457, 4567.47429841396, 4525.29911632283, 
    4491.88683519796, 4438.56575033615, 4376.05347162414, 4397.53773613661, 
    4448.44294110018, 4465.82673511068, 4487.90483830889, 4446.03019810672, 
    4419.18185522252, 4389.95757933208, 4400.61145217698, 4359.28663240238, 
    4227.02127008732, 4009.58021347401, 3850.92644994345, 3640.36848450523, 
    3600.50646255756, 3404.79193203378, 3411.42524954005, 3505.04889666923, 
    3595.30818250343, 3630.04276897278, 3662.87156055393, 3698.45938621674, 
    3757.57710755349, 3813.93134683241, 3853.46858625518, 3842.71186602633, 
    3785.75072588312, 3726.83907291156, 3633.3896253915, 3560.79701475681, 
    3500.59932742814, 3465.77734909714, 3433.39816852821, 3394.10728939141, 
    3337.91649604299, 3264.96653512902, 3227.60742504944, 3218.89441523156, 
    3277.48793660495, 3365.87994586474, 3451.92825462759, 3546.01723933273, 
    3653.69830730641, 3744.70002689153, 3815.57296060554, 3855.0747961651, 
    3882.15136974841, 3917.80105956191, 3944.46627954774, 3974.49122183058, 
    3999.28689295864, 4018.19577927665, 4023.86392130926, 4022.07676969756, 
    4008.52311673209, 4028.26058857903, 3996.7627329067, 3972.4513454536, 
    3979.16388233589, 4021.00105840625, 4081.95658799495, 4121.32121897307, 
    4147.43518521634, 4155.70068090663, 4135.21046129397, 4108.427640587, 
    4035.52513968337, 3911.21130611596, 3619.61370422824, 3389.4954418509, 
    3403.56878860072, 3836.03735074644, 4196.93822408799, 4467.73093852701, 
    4613.73163854618, 4647.00861873546, 4616.34023788518, 4505.88492160577, 
    4521.71031948512, 4299.33848598812, 4323.94658211696, 3576.05189933552, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 1331.292985637, 
    2083.35328286945, 2724.60632207721, 3281.99565932736, 3706.30860675075, 
    3994.1921049613, 4175.74815860626, 4311.35009437805, 4475.63220170032, 
    4668.81594462175, 4900.62590355244, 5089.29154622386, 5222.39184392736, 
    5325.38191624059, 5363.71253583232, 5348.87767104924, 5297.26312656471, 
    5230.48943887263, 5116.20749639511, 4996.88020850463, 4883.65139049892, 
    4742.4110707183, 4575.26971627812, 4398.70021062356, 4225.27744532223, 
    4054.95701387681, 3838.70060363082, 3634.1769090403, 3486.65003141485, 
    3526.46266836441, 3748.89243854119, 4020.03551641621, 4279.28307719042, 
    4519.86174628263, 4702.70676346711, 4825.44395096027, 4940.19303603612, 
    5065.3960872757, 5164.49135605501, 5226.38189949943, 5299.33278370871, 
    5346.753949665, 5325.12530789382, 5178.88343489817, 4865.73496046695, 
    4384.94016791776, 3883.55232282392, 3598.41407577973, 3560.09268641675, 
    3693.24239502579, 3481.60683535961, 2937.72592357591, 2237.34811537208, 
    1447.8666659661, 835.034851901772, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 1199.58146437838, 
    1867.58127540799, 2442.33960108955, 2781.71806018571, 2870.19871331391, 
    2920.3432979712, 2794.52554955815, 2486.99676179934, -0, -0, -0, -0, -0, 
    2983.75445011369, 3900.80046296149, 4369.02598804235, 4693.19659792513, 
    4676.35560830907, 4419.18185522252, 4194.23277779284, 3906.12891061253, 
    3999.64843315678, 4139.64910295478, 4208.7237589253, 4191.48638320263, 
    4150.02206633039, 3997.71656052997, 3841.60682232298, 3700.70618870983, 
    3562.82331206121, 3430.14754148625, 3305.59869916446, 3171.11123979999, 
    3082.19561456491, 3157.52666341367, 3389.89967599493, 3695.92075568186, 
    3932.5603433408, 4097.35439556069, 4191.92514029238, 4293.52641440925, 
    4405.64762145109, 4508.05387791363, 4611.41318207777, 4674.65473653576,
  4819.32791958883, 4847.55730221816, 4877.32792631986, 4761.41850543961, 
    4664.85195658168, 4349.49886116019, 3975.97476324314, 3333, 
    3929.09267354269, 4384.71706056765, 4687.31161391907, 4872.73002476845, 
    4994.02014585344, 5070.70401911108, 5161.91375714763, 5256.09665581671, 
    5406.32505726768, 5500, 5500, 5500, 5500, 5500, 5340.20863548546, 
    5022.15176648433, 4861.91022515031, 4937.44884675988, 4951.89299592686, 
    4873.96119049971, 4749.42758366544, 4562.08649698018, 4164.91531815075, 
    3261.31912627723, 2214.03642479706, 1478.68884277344, 855.295364272955, 
    120, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 100, 170, 
    386.499133726878, 545.419436106388, 1324.25608468959, 1994.71637838929, 
    2550, 2550, 1893.53001652458, 1584.39310898899, 1649.49011671483, 
    1762.93779400443, 1846.00111631343, 2323.87750335617, 2279.05808500641, 
    2279.05808500641, 2174.08020638627, 2353.46705536584, 2363.65495714421, 
    2363.65495714421, 2695.50666974581, 2714.34555090062, 2926.12469139439, 
    3014.24936676646, 3025.10225621468, 3034.34964733199, 3102.65983992087, 
    3117.66286187926, 3264.49932391275, 3187.0835262694, 2877.79165884739, 
    2305.95996082419, 1941.95325919772, 2028.88634049358, 2095.67008549412, 
    2472.68307817313, 3266.92849744038, 5005.658933575, 5409.83324993272, 
    5500, 5483.32364049079, 5363.79010798432, 5349.28191204914, 
    5342.70386114729, 5291.93793147425, 5194.3809349354, 5103.22224646129, 
    4989.89811231253, 4857.93685847825, 4752.7293128579, 4617.33558031335, 
    4508.53533301493, 4525.4748323599, 4495.87587633646, 4516.22890808868, 
    4555.62857972944, 4571.06691859978, 4486.28276507562, 4369.50435350424, 
    4345.37802910977, 4299.29454094438, 4343.71946680647, 4433.32883533073, 
    4444.2211802683, 4423.7130800685, 4368.22596471539, 4325.47915760073, 
    4298.6748137077, 4249.37565214141, 4155.62897744246, 3962.41685958584, 
    3765.41147071606, 3545.47014483236, 3427.83354072401, 3442.89829311604, 
    3557.73568579779, 3594.03413228224, 3643.49570895842, 3683.39377691141, 
    3662.87156055393, 3813.64485742938, 3910.00917345239, 3966.14332641794, 
    3957.13084596345, 3920.61374188302, 3849.776529406, 3789.17664298384, 
    3657.34892267489, 3582.78659957721, 3517.89434496017, 3489.52373819784, 
    3457.22705297292, 3420.13831109361, 3377.15686231386, 3293.4101530799, 
    3245.26902193559, 3210.64882459986, 3255.94372810836, 3340.4846642843, 
    3425.41398737968, 3537.44214759316, 3658.6748098191, 3757.74236614034, 
    3832.40738273374, 3873.41883693442, 3905.00086840166, 3946.68996638148, 
    3989.07774376823, 4023.78023064999, 4047.45800737217, 4073.82811467319, 
    4083.14912962327, 4065.89147763595, 4087.76800013981, 4098.35514623485, 
    4065.89147763595, 4026.54447007219, 4021.11626663601, 4087.07072838132, 
    4136.97175126915, 4180.35297061293, 4218.86824999794, 4229.31081796839, 
    4222.20561884535, 4239.59216349483, 4213.35944123835, 4110.6139657154, 
    3875.9147168786, 3615.92239378233, 2075, 3700.26678232462, 
    4068.13841853297, 4346.82046300842, 4570.48811967065, 4671.81866969785, 
    4716.71022620217, 4640.65484196307, 4634.22335035148, 4321.49713536584, 
    4266.17738799091, 3195.41188711166, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 1065.80177610638, 1798.40011949406, 2377.89260919737, 
    2874.2717244334, 3430.48919278148, 3721.27612304688, 3867.66734233421, 
    4071.54579274883, 4320.71950174819, 4481.7144107472, 4755.15878909484, 
    4905.4699284809, 5102.72217846492, 5260.1826315268, 5341.56974809045, 
    5348.42129348639, 5297.69949740547, 5233.0781243306, 5157.5683092303, 
    5084.23782222658, 4971.59871328779, 4742.4110707183, 4589.96982230177, 
    4356.54764715262, 4217.59519530903, 4048.64329214525, 3850.51198654361, 
    3608.64015041273, 3434.31356095714, 3427.8500105299, 3639.19918959894, 
    3905.82517741705, 4190.53178136803, 4420.20893683752, 4622.56294827644, 
    4800.29532083081, 4940.20402751165, 5046.79269927597, 5143.41858983545, 
    5197.7902416271, 5292.70187551789, 5376.39743053859, 5383.54027740784, 
    5324.32103564432, 5106.01649590208, 4697.55173274604, 4335.33849776841, 
    4077.39112132637, 3737.05313665632, 3480.42376023994, 3189.68072858415, 
    2553.55122375072, 1853.56095484627, 1101.54602050781, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    926.535123984995, 1615.91621584468, 2191.85384798669, 2556.17789953264, 
    2782.94109677749, 2786.24450037171, 2638.28241477722, 2297.51137885108, 
    1659.43101440721, -0, -0, -0, -0, 2536.33867620827, 3752.45595286944, 
    4357.90552560923, 4652.90505455916, 4726.240949108, 4483.05161799804, 
    4160.07235085993, -0, 3829.29732430133, 3748.31139136736, 
    3931.3062225076, 3940.05358055618, 3932.81536592045, 3815.6282833287, 
    3614.5682223014, 3387.2978515625, 3241.02053383166, 3150.80293603859, 
    3065.78548661781, 3000.56346111284, 2997.75167220404, 3181.31401958047, 
    3435.10605237661, 3731.66501335275, 3992.67425354305, 4207.22343761045, 
    4299.1931980505, 4399.7998978106, 4529.03645168398, 4638.65291794403, 
    4718.49837806282, 4779.44385110665,
  4899.8, 4933.9, 4966.4, 4891.7, 4759.3, 4439.6, 4009.3, 3426.9, 3861.3, 
    4360, 4716.8, 4927.7, 4992.3, 5107.1, 5208.3, 5323.1, 5453.2, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5181, 5218.7, 5220, 5131.6, 4959.6, 4670.6, 
    4170.2, 3350.7, 2383.8, 1636.2, 1142.2, 120, 80, 80, 50, 0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 40, 100, 170, 621.7, 712.8, 1608.9, 2169.8, 
    2550, 2550, 2160.5, 90, 2037.5, 2181.4, 2324.1, 2404, 2404, 2595.6, 
    2666.1, 2860.1, 2865.2, 2517.7, 2537.7, 2647.5, 2848.1, 2953.5, 2960.3, 
    2947.2, 2940.6, 2886.9, 2868, 2712.5, 2539.2, 2124.1, 1790.2, 2001, 
    2060.8, 2323.2, 2919.1, 4419.181640625, 5500, 5500, 5307.8, 5109.8, 
    5195.2, 5257.1, 5249.8, 5183.5, 5088.2, 4974, 4846.1, 4783.4, 4665.6, 
    4538, 4522.7, 4506.5, 4530.7, 4553.7, 4537.6, 4438.3, 4289.7, 4128.8, 
    4123.1, 4133.4, 4211, 4230.1, 4290.4, 4235.6, 4166.5, 4110.6, 4053.8, 
    3890, 3733.5, 3510.7, 3481.5, 3434.8, 3424.3, 3508.2, 3561.6, 3672.3, 
    3773.3, 3813.3, 3930.7, 3978.8, 3997.6, 3978.5, 3926.2, 3837.7, 3763.7, 
    3650.3, 3601.9, 3550.1, 3521.3, 3489, 3446.6, 3390.5, 3308.2, 3238.6, 
    3193.2, 3210, 3290.5, 3394.8, 3518.3, 3642.5, 3757.8, 3842.3, 3893.5, 
    3929.4, 3958.41550076125, 4007.10371205604, 4037.3, 4071.1, 4097.3, 
    4115.2, 4115, 4134.1, 4132.6, 4097, 4065.89135742188, 4071.7, 4136.6, 
    4194.7, 4228, 4261.8, 4269.6, 4282.6, 4306.3, 4310.4, 4256.8, 4090.8, 
    3889.6, 3031.5, 3700.26678232462, 3754.1, 4182.9, 4405.1, 4556.7, 4669.9, 
    4636.6, 4516.6, 4233.4, 3968.8, 2709, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 1359.1, 1887.5, 2656, 3316, 3721.3, 3952, 4121.4, 4313.1, 
    4473.8, 4712.2, 4889.9, 5085.4, 5239.6, 5333.2, 5352.7, 5307.5, 5242.6, 
    5151.4, 5051, 4918, 4717.1, 4487.7, 4232.1, 4065.89135742188, 3892.1, 
    3708.8, 3483.7, 3319.5, 3349.8, 3569.9, 3849.6, 4132.5, 4363.1, 4554, 
    4736.8, 4878.6, 4982, 5042.8, 5120.9, 5233.5, 5500, 5406.3, 5500, 5252.1, 
    4996.6, 4740.1, 4509.7, 4201.2, 3840, 3306.1, 2511.2, 1697.125, 170, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 70, 834.803854551359, 1852.2, 2522.95436253561, 
    2688.80567277747, 2688.80567277747, 2638.28241477722, 2250, 1623.9, -0, 
    -0, -0, -0, -0, 3519.8, 4223, 4578.1, 4734, 4585.9, 4334.2, 
    4246.25347954186, 3829.8, 3462, 3565.7, 3609.4, 3687.2, 3626, 3485.8, 
    3255.6, 3118.9, 3015.1, 2988.6, 3019.8, 3099.5, 3312.7, 3582.9, 3868.5, 
    4081.2, 4277.9, 4371.4, 4495.6, 4621.01910701073, 4716.91832585084, 
    4792.2, 4850.3,
  4980.3292459445, 5020.15751938861, 5055.5679085809, 5022.03281946452, 
    4853.79194789034, 4529.76587754787, 4042.60306784274, 3520.88531282084, 
    3793.50805140909, 4335.31315739893, 4746.28108161801, 4982.71910716883, 
    4990.55694303488, 5143.41858983545, 5254.6969385697, 5390.12008034163, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5488.06330471816, 5389.33010022573, 5169.81543941624, 4779.07571895829, 
    4175.50665859157, 3440.1519633162, 2553.62916032264, 1793.6112770465, 
    1429.15591895836, 1122.1259380155, 846.653055803787, 618.596519280046, 
    387.439653279541, 220, 130, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    382.340288811397, 425.785466617812, 495.553629324057, 630.368481982803, 
    856.822549435097, 1280.12060546875, 1893.58970625818, 2344.96349433972, 
    2550, 2550, 2427.56243798484, 2193.79007360743, 2425.52066982558, 
    2599.79107039707, 2802.22419962429, 2790.62281701295, 2529.04103417559, 
    2912.18587715416, 3158.11920992881, 3366.79366386314, 3366.79366386314, 
    2671.78286858751, 2379.92794405606, 2580.64059191887, 2770.12602976525, 
    2892.65803426023, 2895.42332148391, 2860.12506647933, 2778.58573177594, 
    2656.21961486239, 2471.58674475181, 2237.8278442741, 2200.59144226142, 
    1942.24477621766, 1638.44894457643, 1973.17831092378, 2025.90294814803, 
    2173.66380064908, 2571.35767339494, 3815.27745414145, 4922.40904192454, 
    5132.27477086741, 5132.27477086741, 4855.7919319837, 5041.03421752499, 
    5171.46064342578, 5207.58513222988, 5172.70992308385, 5073.09333808727, 
    4958.00549059767, 4834.34046579061, 4814.04319698833, 4713.86000970218, 
    4567.43282397921, 4520.01382495293, 4517.02965998053, 4545.11673789275, 
    4551.72427878011, 4504.20805331895, 4390.34250961319, 4209.89250414037, 
    3912.26727440808, 3946.83934097569, 3922.9854276939, 3988.70983140193, 
    4015.93749454096, 4157.03374963039, 4103.06578848843, 4007.4641410627, 
    3922.56371167985, 3858.13311995435, 3624.39935212604, 3504.51840389404, 
    3255.88926202236, 3417.60548126407, 3441.85892254966, 3405.68848073015, 
    3458.75514593535, 3529.13043550954, 3701.14390947565, 3863.18447882779, 
    3963.74116639532, 4047.67567121536, 4047.67567121536, 4029.15645637134, 
    3999.89640861813, 3931.86770698451, 3825.55766050299, 3738.1842254169, 
    3643.34441077864, 3620.96071875393, 3582.35730256968, 3553.14505730042, 
    3520.71525817508, 3473.08173599618, 3403.87819693304, 3322.97975530361, 
    3231.97273582535, 3175.76853445716, 3164.1465756666, 3240.51223389136, 
    3364.16572711385, 3499.07727531132, 3626.41314841462, 3757.8194050756, 
    3852.12969251304, 3913.6150755017, 3953.76524490166, 3992.71506127885, 
    4029.90401856669, 4050.79752644812, 4094.79424762799, 4120.71581299707, 
    4147.15549342797, 4164.15130860754, 4180.44156961022, 4166.79280243452, 
    4128.08235465518, 4094.62583087218, 4122.22653043781, 4186.17702120252, 
    4252.4261957526, 4275.71653782216, 4304.72821979732, 4309.91711923443, 
    4342.89483041454, 4373.08598819292, 4407.45618460961, 4403.03807956121, 
    4305.71427561558, 4163.22137110477, 3988.06928787908, 3837.94465755304, 
    3440, 4018.99654267093, 4239.79659935068, 4441.67808327036, 
    4623.16936886327, 4632.47972061769, 4398.92782564504, 4145.28450977211, 
    3671.34045720142, 2222.6807040046, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 919.777561694523, 1397.18067919919, 2437.77729879913, 
    3201.51283511651, 3721.27612304688, 4036.24563913452, 4171.30715381099, 
    4305.52515189185, 4465.95014089593, 4669.32082437609, 4874.25707711893, 
    5068.05545173389, 5219.00802010619, 5324.8158023114, 5357.00249959007, 
    5317.22298437148, 5252.20002359477, 5145.22849959196, 5017.66457535914, 
    4864.38201937079, 4655.08477099385, 4385.3385316582, 4107.71519192101, 
    3910.6876526659, 3735.47306075624, 3567.09603730106, 3358.74913596743, 
    3204.69155246331, 3271.77326246576, 3500.52164408084, 3793.3088022128, 
    4074.53579172404, 4305.90590717307, 4485.51084149148, 4673.28059322413, 
    4816.99019742938, 4917.12867887675, 4942.26089937211, 5043.99788505255, 
    5174.38465338656, 5316.94067687406, 5429.05204926276, 5462.49308876518, 
    5398.25732065627, 5295.55997169833, 5144.76336082456, 4941.98908354189, 
    4665.43898307603, 4199.54409773268, 3422.54177224637, 2468.77357721399, 
    1537.41766014626, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 834.803854551359, 
    1512.50279851896, 2005.83190586972, 2309.44840269853, 2450.54710920634, 
    2250, 2250, 1588.28199275357, -0, -0, -0, -0, -0, 3287.09259127595, 
    4088.03424409215, 4503.30076826239, 4741.68777585758, 4688.77648167513, 
    4508.33631284944, 4163.42869833995, 3830.2164120184, 3175.73134948332, 
    3200.12990189844, 3278.69814146574, 3441.58611327241, 3436.44920966913, 
    3357.00244385341, 3123.98828960563, 2996.81560086289, 2879.42489171357, 
    2911.39004545303, 3038.96099508715, 3201.28668168151, 3444.0152699223, 
    3730.69905054341, 4005.27627944144, 4169.75298944188, 4348.54152419149, 
    4443.52721749509, 4591.44481763477, 4685.33696237877, 4779.07571895829, 
    4865.94993953278, 4921.07834480866,
  5032.92867588349, 5085.99160682556, 5126.99764012024, 5118.25185268652, 
    4955.03149826151, 4612.25422965695, 4149.79003773736, 3666.57843477256, 
    3798.61240153853, 4386.49768838833, 4790.73295568097, 5074.77398404932, 
    5101.07760722581, 5151.59502970023, 5336.10084179103, 5448.00507575219, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5357.1985024792, 5069.73360697899, 4553.73572169029, 3946.89973011609, 
    3116.81600753047, 1907.46006121315, 1907.46006121315, 1750.31019740495, 
    1512.82691561821, 1208.94199835615, 738.619525162333, 220, 130, 120, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 150, 603.300191235082, 667.508531967295, 
    538.200910062152, 630.368481982803, 856.822549435097, 1405.68699995804, 
    2089.78778032001, 2418.49920202865, 2550, 2622.83553886791, 
    2747.8089361534, 2773.53299769021, 3040.80368594565, 3091.59270903075, 
    3158.06599430688, 3120.65220112486, 3046.57012854129, 3300.45336759044, 
    3550.99061943318, 3612.57227319316, 3366.79366386314, 2583.36356655798, 
    2400.82000321383, 2552.11898268036, 2784.06999975711, 2907.62893445192, 
    2871.6020148564, 2791.22940050275, 2617.83090930657, 2406.9087257915, 
    2054.27696907627, 1827.45701699937, 1802.07722478058, 1683.16320530693, 
    1638.44894457643, 1982.53047739804, 2052.58233396938, 2173.66380064908, 
    2466.66776221529, 3387.2978515625, 4570.67400169003, 4929.17701617885, 
    5039.6316840347, 4874.05659929983, 5003.20662467964, 5190.70542015141, 
    5254.56948305078, 5233.42877513996, 5091.03880916715, 4946.43218540326, 
    4869.48141225681, 4855.87764458452, 4741.41730559854, 4741.41730559854, 
    4677.9580673091, 4602.66855499778, 4572.15342275341, 4548.75240986906, 
    4406.50049792499, 4210.90639867467, 3996.61253584561, 3878.25945314569, 
    3768.84887351141, 3686.0522931149, 3790.89992786817, 3881.22542635781, 
    3834.83808676935, 3723.29919434665, 3575.43628080012, 3503.35314493835, 
    3362.53579835637, 3264.43594774861, 3190.87526220851, 3269.0106992718, 
    3255.88926202236, 3335.32658255232, 3358.08377269987, 3633.63275177696, 
    3772.9613657307, 3900.19733732051, 4017.90396174952, 4076.09771307239, 
    4094.19027030455, 4080.22089113606, 4038.29626475461, 3974.42530039383, 
    3889.38433568047, 3794.89760274705, 3735.86531051537, 3672.46369138211, 
    3633.36624065702, 3606.42788759536, 3584.7787872093, 3542.25834512845, 
    3479.05288029687, 3391.22777570153, 3303.02173649156, 3208.28202420204, 
    3141.95007949751, 3127.86391394516, 3201.89154583324, 3321.77767865535, 
    3468.18679321538, 3612.40977071374, 3747.37031016194, 3841.4289419057, 
    3903.73995636773, 3958.35467933246, 3988.8221549478, 4017.91902147464, 
    4045.04651340067, 4065.89147763595, 4085.04570218883, 4109.17367020303, 
    4127.8831556665, 4145.10830176833, 4138.81070296011, 4115.68239757757, 
    4077.38055957312, 4150.52405706573, 4222.70115792022, 4295.42324276613, 
    4323.25078427377, 4340.02160638574, 4360.08916766444, 4388.22923345963, 
    4419.47427712142, 4456.5531290085, 4479.87046529089, 4455.38677328812, 
    4365.83591211795, 4210.93697663841, 4031.98868372499, 3440, 
    3855.44378345404, 4047.89253235506, 4271.40629722256, 4397.50853751434, 
    4397.50853751434, 4293.27688806588, 3998.44703920921, 3001.21919635974, 
    2222.6807040046, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    803.625015916513, 1322.4191623767, 2282.6117565196, 3138.47357284546, 
    3743.6267201192, 4126.20372490787, 4296.75775721215, 4438.55149227736, 
    4570.04356473396, 4722.90301398617, 4914.10141306441, 5094.92651030501, 
    5244.87731201616, 5353.05291515663, 5375.84810952719, 5325.02563145418, 
    5223.88292589973, 5052.58733139336, 4906.88565386762, 4753.08678812208, 
    4541.95514325494, 4257.2064976903, 3972.07244786874, 3745.90169608509, 
    3563.829470016, 3419.29985654414, 3281.63049508576, 3160.54182277081, 
    3301.18429917327, 3513.09743538677, 3748.80994096388, 3974.95094852771, 
    4188.00713874299, 4382.28746143231, 4588.52246421888, 4749.34922952819, 
    4871.03011150962, 4923.19668346307, 5010.92809113102, 5147.74850582385, 
    5325.62869870416, 5445.44727677905, 5500, 5483.4555306875, 
    5428.46371307143, 5346.35417723749, 5178.29041440167, 4873.78506705715, 
    4406.05028682184, 3689.86845933493, 2900.14293937558, 1537.41766014626, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 1222.92144943369, 1790.1895439141, 
    2119.4774096446, 2119.4774096446, 2250, 2250, 1445.5815868833, -0, -0, 
    -0, -0, -0, 2948.94993712953, 3906.47651775969, 4356.91661523523, 
    4645.43161237684, 4712.12506917661, 4580.24572181732, 4309.77726942309, 
    3928.61362584876, 3407.06152881074, 2982.26182794897, 2930.80898280466, 
    3190.00725508879, 3292.72764214919, 3354.84232654471, 3300.23253893122, 
    3140.66439292298, 2998.91744332321, 3002.68153516178, 3105.42384728962, 
    3313.6860923149, 3629.53986665854, 3915.85697769617, 4151.29839259132, 
    4324.53002107108, 4473.18007927199, 4574.26378068077, 4644.17036947649, 
    4732.29382088274, 4811.80284639711, 4893.131673557, 4952.4686335588,
  5044.8, 5098.8, 5119.3, 5098.2, 4936.6, 4561.5, 4092.3, 3640.4, 3749, 
    4419.4, 4830.1, 5110.1, 5143.41845703125, 5206.9, 5314.9, 5500, 5500, 
    5493.5, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5428.6, 5500, 4876.5, 4335.1, 3599, 2719.7, 2695.7, 2662.3, 2517.9, 
    2225.7, 1539.6, 50, 120, 120, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 0, -0, -0, -0, -0, -0, -0, 150, 833.7, 845.9, 
    853.6, 854.2, 955.6, 1808.7, 2412.2, 2702.3, 2760.8, 2789.1, 2886.7, 
    2998.8, 3262.9, 3445, 3557.4, 3524.9, 3480.6, 3622.7, 3685.4, 3570, 
    3085.4, 2503.1, 2534, 2697.5, 2898.4, 2948, 2881.6, 2790.5, 2611.1, 
    2370.56158557313, -0, 160, 1025.21479783781, 1583.9, 1697.125, 1974.1, 
    2107.96239883132, 2107.96239883132, 2494.2, 3200.3, 4383.1, 4804.2, 
    4945.4, 4932, 5031.8, 5237.5, 5317.2, 5304, 5500, 5081.2, 4953.9, 4900.6, 
    4848, 4848, 4782.4, 4705.4, 4610.8, 4508.1, 4329.6, 4180, 3967.9, 3769.6, 
    3721.27612304688, 3647.6, 3659.3, 3576.3, 3348.3, 3019, 3002.4, 3001.3, 
    2986.4, 3000.3, 3001.5, 3112.4, 3241.8, 3455, 3612.5, 3834.9, 3949.5, 
    4033.5, 4084.2, 4101.7, 4088.5, 4065.89135742188, 4008.3, 3938, 3856.4, 
    3773.1, 3728.6, 3681.5, 3643.9, 3615.6, 3577.8, 3539.3, 3482.8, 3398, 
    3310.2, 3217.4, 3144.1, 3119.8, 3183.2, 3307.2, 3453.8, 3593.5, 
    3721.27612304688, 3797.7, 3863.2, 3910, 3953.9, 3979.8, 3992.6, 3977.5, 
    3981.1, 3991.2, 4006.5, 4034.4, 4035.1, 4047.1, 4053.4, 4135.1, 4212.5, 
    4283.3, 4328, 4349, 4372, 4406.3, 4455.1, 4509.6, 4548, 4540.6, 4488.3, 
    4362, 4188, 3768.5, 3836.5, 3836.8, 4004, 4195, 4218.6, 3908.9, 
    1896.03911720189, 70, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 1587.7, 2528.8, 3306.7, 3888.9, 4223, 4381, 4517.6, 4650, 4799.7, 
    4967.3, 5143.41858983545, 5281.1, 5371.9, 5377.3, 5295.8, 5183.7, 5005.5, 
    4866, 4710.8, 4494.3, 4218.1, 3935.9, 3693.9, 3495.3, 3326, 3225.5, 
    3193.7, 3326.4, 3530.2, 3740.3, 3932.4, 4108.4, 4287.3, 4485.1, 4677.9, 
    4836.1, 4928.4, 5044.4, 5174.2, 5339.9, 5500, 5500, 5500, 5500, 5500, 
    5215.8, 4932.6, 4500.8, 3823.5, 3065.78540039062, 1059, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 40, 565.376620444443, 1958.5541560972, 2119.44993275496, 
    2250, 2250, 1250, -0, -0, -0, -0, -0, -0, 3551, 4192, 4503, 4647.4, 
    4568.7, 4365.2, 4037.2, 3540.6, 2980.7, 1902, 2768, 3065.8, 3295.2, 
    3295.2, 3266.1, 3117.7, 3078.8, 3163.7, 3387.2978515625, 
    3721.27612304688, 4023.6, 4285.2, 4466.7, 4600, 4681.9, 4742.6, 4803.9, 
    4848.1, 4912.1, 4973.6,
  5056.76932243833, 5111.54618039021, 5111.54618039021, 5078.24749503872, 
    4918.25744326612, 4510.80454026882, 4034.76654302428, 3614.19063912455, 
    3699.48550928694, 4452.25249926604, 4869.56031715392, 5110.1, 
    5173.9963142228, 5262.2173786553, 5293.7929397493, 5430.91332787923, 
    5425.09044654863, 5486.91116876777, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5421.39257776028, 5199.31596118267, 
    4723.21021245647, 4081.15112967156, 3531.96023692031, 3483.9081215267, 
    3574.21785786591, 3522.90320273947, 3242.45307021751, 2340.60044576711, 
    1422.07186637295, 806.226855052668, 388.589231969222, 220, 90, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 60, 60, 60, -0, -0, -0, 
    -0, -0, 1065.13999018601, 1064.02640010958, 1024.36768255671, 
    1049.01333931092, 1258.09536998652, 1646.38481505787, 2211.63703163277, 
    2734.57596636045, 2986.0794993596, 2971.58676265889, 2955.36382697119, 
    3025.62532076787, 3224.12947072977, 3485.01385375916, 3798.36368196785, 
    3956.69610419615, 3929.07928363366, 3914.67964350191, 3945.01755772368, 
    3622.7, 3527.34743282107, 2782.04296263851, 2422.81360052491, 
    2667.17369501951, 2842.87362696265, 3012.73528672141, 2988.34664131686, 
    2891.53469443837, 2789.70951314374, 2604.43714048112, 2334.20749278165, 
    1898.44211827902, 1542.58715923581, -0, 1484.68816907211, 
    1740.72116017347, 1965.60894138933, 2107.96239883132, 2147.5339468221, 
    2521.68042209255, 3013.25678062404, 4195.61897271538, 4679.15836122614, 
    4851.133867915, 4989.98803355365, 5060.40211212047, 5284.33790487616, 
    5379.8544139237, 5374.53682001959, 5330.85808027182, 5216.05781904441, 
    5038.28666994432, 4945.27459829145, 4954.53805110375, 4954.56042926009, 
    4886.93878440509, 4808.05749106325, 4649.39481348018, 4467.48573117766, 
    4252.61311231703, 4149.10584682841, 3939.14882796382, 3660.92726889355, 
    3660.92726889355, 3609.10911843915, 3527.6298026413, 3271.34685861746, 
    2861.8031156689, 2314.63424913702, 2429.29801285032, 2499.20868368662, 
    2610.31683337247, 2736.07304259679, 2812.07213423353, 2955.83641248066, 
    3227.64420082699, 3574.62512040964, 3866.95972731319, 4036.24926333881, 
    4126.13528390447, 4166.82343836524, 4150.44929999598, 4127.40039996778, 
    4082.89946671572, 4033.01890943504, 3978.32145364795, 3901.52347547208, 
    3823.44449444591, 3751.27679825902, 3721.27612304688, 3690.44708675532, 
    3654.34262412183, 3624.70596345738, 3570.88709966655, 3536.28169450036, 
    3486.6142577909, 3404.72373781175, 3317.35138922102, 3226.422589815, 
    3146.33989789732, 3111.67146228262, 3164.49101983856, 3292.67553629151, 
    3439.4531716411, 3574.49286648566, 3685.36600839485, 3753.9560393101, 
    3822.74742221282, 3861.67618242377, 3918.89068000554, 3941.76250893052, 
    3940.21175951028, 3889.19635746434, 3877.05795970386, 3873.24998849618, 
    3885.21074866886, 3923.77865196509, 3931.46343198121, 3978.47631874437, 
    4029.46547321509, 4119.58299228302, 4202.33015022304, 4271.11779831345, 
    4332.83141017334, 4357.92347112883, 4383.86896305177, 4424.43865590767, 
    4490.77399004562, 4562.60099478045, 4616.035222974, 4625.79268909784, 
    4610.79732273264, 4513.00247007362, 4343.91243405158, 4096.9678572344, 
    3817.64294477621, 3625.72143804519, 3736.60372953589, 3992.44584946079, 
    4039.62373853847, 3524.58414949955, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 1852.93187624811, 2774.97022424922, 
    3474.99723774056, 4034.19110822047, 4319.73764273154, 4465.32714308645, 
    4596.71613126888, 4730.01646861658, 4876.42529288602, 5020.40364951388, 
    5187.72584539554, 5317.35768943021, 5390.70754526109, 5378.68214902704, 
    5266.62852834647, 5143.41858983545, 4958.37407797266, 4825.12380894111, 
    4668.46830199904, 4446.67809151248, 4179.08714972309, 3899.6661237447, 
    3641.85519254873, 3426.80484466673, 3232.75638498102, 3169.2764013265, 
    3226.76533612161, 3351.55277887041, 3547.33468445097, 3731.73379284763, 
    3889.7867954879, 4028.80674855647, 4192.23927068536, 4381.59166730582, 
    4606.42910709273, 4801.10687164601, 4933.57460412379, 5077.79201429083, 
    5200.6701883743, 5354.2674465104, 5464.65866686568, 5500, 5500, 5500, 
    5412.04248344969, 5253.35350900251, 4991.37690046479, 4595.64250486362, 
    3957.19884970778, 3217.63013097644, 2180.60948245598, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 1964.12344621424, 2250, 2250, 1679.38359590569, 
    1463.64291582816, -0, -0, -0, -0, -0, 3195.58964421974, 4027.15257766301, 
    4360.62090611149, 4582.74959056834, 4557.05732670339, 4392.56003508355, 
    4145.8370305113, 3674.17989324933, 2979.11959495284, 2073.20665780415, 
    2345.96072348596, 2838.9356807289, 3235.50961338387, 3461.49904562595, 
    3391.59122419243, 3236.38468048116, 3154.9943442454, 3222.04527923043, 
    3453.36253506423, 3810.12749885282, 4131.33557382584, 4419.18185522252, 
    4608.82342106985, 4726.89849941386, 4789.51560706108, 4841.04906254948, 
    4875.41408467523, 4884.44446435777, 4931.03432956596, 4994.79532997288,
  5023.44759176876, 5026.29963171568, 5118.11090407112, 4979.36262911642, 
    4791.36597504497, 4444.75033377513, 3989.38246714818, 3434.86393432836, 
    3560.75949444583, 4585.69152438164, 4945.62857743526, 5097.65475409155, 
    5097.65475409155, 5292.65650916622, 5242.4296131648, 5398.79306784713, 
    5292.76529429391, 5379.8570449381, 5468.66888810767, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5475.84726644584, 5425.41412739273, 
    5331.20238233828, 4914.30013919355, 4290.7638740685, 4055.28862534487, 
    4483.68817394872, 4677.56740640126, 4658.76326975034, 4390.30063697468, 
    3459.79680407309, 2058.6967413833, 1111.38285130325, 526.600413818677, 
    306.080280434948, 110, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 50, 70, 80, 80, 60, -0, -0, -0, -0, 1467.86743231721, 
    1335.79139062099, 1344.5345522559, 1348.49393071173, 1659.87386652379, 
    2046.14284683438, 2790.37366250889, 3408.58419780517, 3505.42292836256, 
    3303.55910512292, 3094.23316688248, 3023.04520253836, 3287.49319798829, 
    3478.99691600387, 3849.81367612732, 3965.95144552564, 3965.95144552564, 
    3914.67964350191, 3787.90505840843, 3573.00915078254, 3142.98019328473, 
    2256.09350466087, 2472.25859325978, 2805.36407591694, 3050.75945061425, 
    3166.49099001934, 3085.08477694035, 2942.21326256146, 2867.85625991729, 
    2693.85340885916, 2470.88844964773, 2281.6326416959, 1935.05359591651, 
    1659.12025424165, 1542.64606765131, 1995.47738366991, 2070.11074751043, 
    2173.82011852351, 2234.16818094781, 2524.42031287892, 2785.2916637513, 
    4202.09257172564, 4635.37263913453, 4748.72303269017, 4955.53617496533, 
    5065.13840384699, 5300.78611908347, 5375.43315174839, 5421.56519049176, 
    5372.68887353244, 5276.54498720499, 5081.48574971099, 4892.01026738555, 
    4959.63670770955, 4999.29670319072, 4933.96778971594, 4849.87692123013, 
    4646.79881421256, 4521.35081001848, 4222.53727229091, 4260.78531281206, 
    4176.95321275495, 3920.39550129076, 3881.95332500466, 3769.14396878804, 
    3454.18343894503, 2966.86934426042, 2275.2625933428, 2199.19522704451, 
    2372.68532999417, 2644.34681199945, 2473.70972003787, 2581.85330394111, 
    2593.21633472054, 2987.2460991658, 3461.06724041916, 3810.00632124423, 
    4087.7605798237, 4191.46262551729, 4215.38422468759, 4207.07264276182, 
    4161.24656167294, 4102.74362850074, 4029.66835713951, 3980.98217810988, 
    3967.68157552298, 3890.57540958726, 3813.00416774527, 3726.92410367372, 
    3735.24059826463, 3709.89523072902, 3685.37896532559, 3649.06115555611, 
    3605.58606013839, 3597.30265437909, 3517.16411270728, 3410.67007144892, 
    3318.01393038643, 3228.75338640802, 3140.31835817273, 3113.11823279931, 
    3148.8180319624, 3280.93609123358, 3413.81063422413, 3552.39779191221, 
    3657.28180323434, 3721.27612304688, 3796.2457041992, 3830.02512975096, 
    3941.47489943026, 3951.88054627913, 3855.00744140117, 3797.71646495009, 
    3762.2787246733, 3725.32689300785, 3722.84096599148, 3765.67650683665, 
    3754.04293210683, 3859.06889925437, 3940.28367593748, 4038.37745831453, 
    4153.60192600493, 4224.37596474985, 4289.61988762713, 4324.80078078477, 
    4357.90194641309, 4430.53250528383, 4498.15341811907, 4621.13816447479, 
    4690.34968312288, 4697.60835946642, 4680.42096027205, 4608.33782410329, 
    4481.43745114844, 4289.7553437471, 3887.51908389728, 3437.95150856571, 
    3468.61722592103, 3468.61722592103, 2866.85850361514, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 1755.20850870698, 
    3201.44439063088, 3754.96503992699, 4175.92872581661, 4373.79152744747, 
    4537.11398531201, 4643.8086506879, 4742.34434868894, 4905.82192657106, 
    5055.63414376882, 5220.95980141478, 5340.1805258634, 5441.93068009299, 
    5400.25874000741, 5257.0432450363, 5143.41858983545, 4971.59646447218, 
    4844.54552118867, 4709.4160365354, 4470.57188464448, 4235.95213374914, 
    3951.18461585411, 3678.18140249102, 3431.70848160509, 3235.1213082687, 
    3073.2864887874, 3246.35025586165, 3351.55277887041, 3554.45114037532, 
    3722.32327409228, 3847.15135658557, 4033.28417055992, 4114.26401080236, 
    4071.72422279108, 4560.85220334709, 4793.99203365596, 4940.75402461733, 
    5072.00910907258, 5254.7567845022, 5348.76517782296, 5470.02437781455, 
    5494.1384628282, 5500, 5485.55481058879, 5401.15253099783, 
    5249.36025653842, 4991.34290861954, 4605.13257208691, 4033.83016943915, 
    3371.53284117356, 2180.60948245598, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 1654.53097764754, 2250, 2250, 2214.70019486091, 1613.94917346897, 
    1337.91216635998, -0, -0, -0, -0, 2647.50948429989, 3952.50063154824, 
    4300.8116488482, 4392.56003508355, 4392.56003508355, 4392.56003508355, 
    4260.58590320375, 3832.81497488469, 3089.24972499671, 2073.20665780415, 
    1867.13348438516, 2569.34336542643, 3172.43632438377, 3527.75741167485, 
    3408.6049080465, 3269.89346738251, 3177.70201721436, 3217.76739917073, 
    3453.11195902483, 3796.82026206773, 4128.96190537479, 4469.08999097903, 
    4706.19060065055, 4838.08814666193, 4893.70014113024, 4928.97847489516, 
    4998.28679077241, 4971.27236337062, 4997.16790775416, 4992.99126849293,
  4999.75035993491, 4977.75252329, 4961.83023527355, 4843.33150497072, 
    4590.42029442578, 4171.92809354916, 3589.32942293124, 3436.37207855272, 
    3679.84682069288, 4435.68811887878, 4849.93989805779, 5208.8186890009, 
    5258.28336904514, 5306.27151809559, 5252.9120062607, 5143.41858983545, 
    5148.54468334471, 5208.67499250796, 5384.86719406715, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5441.4842214491, 5309.24186621124, 
    5291.87272464514, 5220.01488986484, 4985.58759385503, 4676.36743990492, 
    4624.10119091841, 4819.97975684739, 5083.14046428388, 5083.14046428388, 
    4819.0245680368, 4035.61140817592, 2777.47187519646, 1669.98996519101, 
    847.170244538767, 434.775341167201, 210, 90, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 0, 50, 60, 70, 80, 80, 80, -0, -0, -0, 1444.88033423125, 
    1760.90699276349, 1737.03484616119, 1879.02895013422, 2116.33021009906, 
    2524.16658770782, 3065.78548661781, 3546.47503692894, 3772.61913655597, 
    3721.27612304688, 3356.60417383112, 3215.59974202433, 3115.50537494283, 
    3160.88599508885, 3373.43632017055, 3617.60224421601, 3965.95144552564, 
    3965.95144552564, 3906.51273877535, 3721.27612304688, 3413.08228549233, 
    2801.79250038168, 2341.02329537218, 2644.5629146365, 2867.9761822337, 
    3117.79045133809, 3174.54954816305, 3098.84128031878, 2990.68463599408, 
    2899.6591226589, 2785.98120462316, 2606.15674803317, 2402.52283103913, 
    2214.75231487212, 2070.48625688001, 2038.29622669264, 2053.31782443073, 
    2085.90514273903, 2288.3561161808, 2469.68623803548, 2822.98024443061, 
    3363.25251353587, 4107.24655446267, 4318.36866383338, 4518.90192961999, 
    4779.07571895829, 4999.1017225057, 5200.19535116557, 5349.21304711937, 
    5426.77934681307, 5333.16183811469, 5123.44850354948, 4909.0147396458, 
    4800.91824677179, 4892.45723173982, 4991.2948041905, 4990.53720052921, 
    4883.46073167794, 4779.07571895829, 4666.91675102261, 4570.89809885142, 
    4462.71946262199, 4388.18249737072, 4217.02904262119, 4002.61188260394, 
    3733.57767669977, 3229.34152438879, 2809.14119649546, 2636.74383516171, 
    2650.21501713571, 2805.87197827273, 3052.28992126699, 3041.96095166038, 
    2953.38410408298, 3036.3741087881, 3314.94913429572, 3659.34131417311, 
    3943.02842845719, 4142.94259129335, 4224.10026836945, 4239.41226348462, 
    4199.99016248308, 4128.74742364884, 4065.89147763595, 4005.43865289481, 
    3987.87600734208, 3953.4506097987, 3894.82618017144, 3819.85890038191, 
    3782.4732771283, 3752.80354291447, 3736.33092806639, 3702.5266019141, 
    3649.66221849325, 3609.33895314673, 3569.46469083131, 3506.01657000486, 
    3410.72268947975, 3311.80119075815, 3225.83467674788, 3150.57569806169, 
    3119.10073689802, 3136.69023581363, 3240.46532782163, 3363.9411730526, 
    3479.13967370885, 3584.41582471272, 3665.89170783764, 3755.61384356662, 
    3848.62123841982, 3915.44120241943, 3972.15400048486, 3948.95241546235, 
    3876.24415378699, 3800.65222875279, 3737.57863531017, 3688.50003382422, 
    3660.46944822574, 3710.38369996553, 3778.96202397539, 3859.44591922391, 
    3951.52404361542, 4044.71930611424, 4114.87459209827, 4171.77092592322, 
    4230.65866524518, 4309.34051442587, 4401.35856325558, 4517.51041147955, 
    4626.32824264881, 4714.49727735702, 4752.36219940783, 4746.62088827757, 
    4682.62680883805, 4566.81420310192, 4366.67157985086, 3961.22794575381, 
    3591.51753950595, 3387.2978515625, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 2466.96645827504, 
    3307.2463988923, 3842.03894205417, 4271.37159416048, 4451.29876055156, 
    4542.52038944936, 4641.33658571009, 4779.07571895829, 4948.25009462553, 
    5114.40700530733, 5244.92639494708, 5327.01341236635, 5373.48538705147, 
    5343.75466593084, 5267.05239691946, 5163.56795854906, 5042.51576482595, 
    4918.60137614713, 4758.50623984568, 4540.0062308613, 4288.84861073454, 
    4012.57261042614, 3731.81727796038, 3444.10319065891, 3220.03851628382, 
    3066.25957982226, 3182.94241584005, 3348.75571509583, 3521.59244998102, 
    3697.3715818192, 3819.16211428228, 3964.57748613689, 4047.2902669779, 
    4217.01153406842, 4466.48968698246, 4733.22933252745, 4935.7163028567, 
    5092.22228244663, 5261.23116332192, 5391.42352338127, 5466.29930332233, 
    5500, 5500, 5479.8956594759, 5387.76270976636, 5209.42267991773, 
    4954.71557227542, 4556.72857964517, 3984.00902676083, 3422.22321775697, 
    2686.12276940066, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 570, 2250, 2250, 
    2665.73242264786, 2550.82377029924, 2342.8063252063, 1939.98080537621, 
    -0, -0, -0, 2659.50859876243, 3785.79690610185, 4244.31033612193, 
    4392.56003508355, 4392.56003508355, 4361.73866084916, 4235.7551182198, 
    3915.57420029477, 3340.93872519992, 2723.99973167114, 1867.13348438516, 
    2466.66776221529, 3081.56376530828, 3412.39778400847, 3430.03588824373, 
    3257.36939487379, 3144.91002882881, 3216.6063142238, 3497.15184113519, 
    3775.56915442706, 4108.41035323455, 4432.19252673438, 4739.62160938982, 
    4914.94577550785, 5009.00669698773, 5041.17098302688, 5053.62043013305, 
    5075.41900622962, 5050.67726123394, 5017.51346004864,
  4965.49508815292, 4948.65074697299, 4899.32275919064, 4747.43512029173, 
    4568.3353361913, 4047.19431689313, 3322.39391693595, 2450, 
    3387.2978515625, 4657.27106789675, 4908.09854425488, 5286.63483435272, 
    5361.9413509289, 5232.7037865541, 5299.51049970051, 4972.46022557423, 
    4968.10359138417, 4930.77579726304, 5319.96194320695, 5493.37718100435, 
    5500, 5240.37128454655, 5312.79938536759, 5500, 5500, 5500, 
    5445.74754129598, 5357.70140725034, 4895.94694139865, 5083.89391933342, 
    5083.89391933342, 5101.01070568268, 4709.36215931821, 4441.04937215467, 
    5087.78981072552, 5419.61150543159, 5495.73822619705, 5287.71007148889, 
    4704.53050170492, 3305.62248194437, 2077.33944384883, 1138.05341922269, 
    508.457852729989, 253.361404418945, 90, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 0, 50, 60, 70, 80, 80, 80, -0, -0, -0, 1565.11631009849, 
    2062.10571047806, 2002.2856765507, 2403.44558392371, 3065.78548661781, 
    3597.28552023755, 3937.85517225735, 3947.30668182314, 3947.30668182314, 
    3956.63787376714, 3230.04343093795, 3263.09908681427, 3314.4183305478, 
    2921.86395554905, 3065.78548661781, 3351.62511415084, 3794.23258247722, 
    3949.72207179109, 3884.32287307431, 3772.11711282765, 3071.54089382072, 
    2763.55067271992, 2341.02329537218, 2691.23206497914, 3037.81933338552, 
    3158.43849851779, 3108.56499986904, 3100.59589804514, 2975.84110107343, 
    2901.93818895269, 2854.00123476002, 2742.9079461097, 2510.24722469092, 
    2313.75717577645, 2181.50493320786, 2169.0120143804, 2139.12840839491, 
    2073.51134657684, 2350.80555342209, 2854.72247948556, 3280.19616889717, 
    3730.766629041, 4082.92675401774, 4065.89147763595, 3986.615886247, 
    4291.1728253929, 4895.92068551698, 5208.8757450648, 5369.20021708155, 
    5379.58423582185, 5280.0784595368, 5020.94093139477, 4537.267848552, 
    4626.36753872213, 4855.65680391184, 4984.02962978081, 5022.564116313, 
    4944.91550350058, 4891.61748198899, 4870.0235009824, 4790.51482747682, 
    4746.99117556287, 4622.3084480904, 4401.02034761284, 4042.49342985201, 
    3730.80876249988, 3393.02940619975, 3105.98658279541, 2969.15529830998, 
    2926.41976154331, 3135.93024623228, 3487.69518057092, 3627.92554566349, 
    3419.48240135322, 3353.20457822831, 3611.40265269949, 3881.88320150579, 
    4067.06556688915, 4199.19279708887, 4264.11179488083, 4247.21780553788, 
    4178.99223694035, 4096.16528293304, 4036.34186200065, 3988.53212502862, 
    3994.0389827649, 3946.96651476178, 3904.78068551345, 3850.29495774303, 
    3808.41979453151, 3767.97507397183, 3742.68584402531, 3693.19280762797, 
    3643.57546499648, 3621.42801935842, 3597.56981324624, 3506.87482594289, 
    3415.44571195962, 3308.38140443181, 3221.14102445776, 3150.99001944991, 
    3100.35072697736, 3090.8064458714, 3206.77424567629, 3313.7598691647, 
    3414.54784622419, 3551.22593711234, 3580.11324332941, 3724.86353442399, 
    3840.28607023162, 3922.00204989032, 4038.80651535454, 4039.3212276793, 
    3955.18913143275, 3867.33918295819, 3779.46858863423, 3694.26064040175, 
    3596.6758542738, 3684.64245924606, 3721.27612304688, 3768.6846332789, 
    3863.40921548702, 3929.16881585707, 4002.7798157068, 4065.89147763595, 
    4150.49680477999, 4229.93013253198, 4374.944066595, 4526.87436223691, 
    4641.84916022221, 4745.24276524702, 4752.59413281134, 4752.59413281134, 
    4752.89816493226, 4669.2715554251, 4366.67157985086, 4022.39928429718, 
    3591.51753950595, 2567.01380318975, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 2466.66776221529, 
    3344.89127701425, 3925.91759373948, 4359.18761426932, 4490.58909897334, 
    4542.71731142236, 4501.24442084582, 4794.53143913104, 4983.71309505579, 
    5163.80670366826, 5258.34760340813, 5298.94798066017, 5363.6007883418, 
    5345.55894163551, 5315.43366774963, 5250.38808866631, 5086.99012159765, 
    4962.07970038704, 4779.07571895829, 4618.09092364133, 4351.06222927534, 
    4098.2591768067, 3815.90810339831, 3480.0932258963, 3162.83368524667, 
    2997.2747360902, 3202.34020339475, 3328.3370797481, 3491.73859517096, 
    3673.84899935564, 3841.08649999383, 3968.64664792385, 4017.35610577739, 
    4124.28223520102, 4424.82223505885, 4700.7546774604, 4882.95853953189, 
    5103.79768699509, 5286.7070599366, 5394.07277996116, 5482.13013984789, 
    5500, 5500, 5483.9953068134, 5399.96969859243, 5208.54966741361, 
    4932.45645481478, 4563.90187602162, 4042.66865189473, 3479.84773570119, 
    2855.7696638481, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 775, 2250, 2250, 
    2967.39726830198, 3002.07577869022, 2844.64996142735, 2406.22743487596, 
    1320.88817369508, -0, -0, 2659.50859876243, 3841.32812654138, 
    4310.73215311716, 4373.33719205212, 4373.33719205212, 4330.08852486073, 
    4256.58368679229, 4051.13761075869, 3642.27420298549, 3140.09731748284, 
    1790.40496324359, 2531.74040679168, 3204.63195544888, 3372.47664161479, 
    3372.47664161479, 3207.05804679099, 2987.94363628477, 3246.35844819827, 
    3483.24648230707, 3783.50990715709, 4080.74157093335, 4394.52274969998, 
    4739.77846196963, 4948.41939594418, 5076.47660180378, 5128.98599533774, 
    5128.98599533774, 5128.98599533774, 5085.03949053607, 5024.94445345409,
  4975.66255769623, 4914.66859118526, 4814.42030956456, 4687.01068896295, 
    4590.60723421944, 4354.14499725315, 3994.78844018355, 3836.30265346653, 
    3501.57949779877, 4449.84393112404, 4852.16476003605, 5232.69943474924, 
    5332.74664037034, 5283.90827933358, 5182.89991758845, 4878.6657375749, 
    4759.33421886516, 4901.28482977121, 5192.63750300709, 5345.46637328909, 
    5365.08910899293, 5143.41858983545, 5088.21726504709, 5214.9989015279, 
    5354.01168702949, 5306.34446156065, 5233.89669242279, 5096.52358219051, 
    4787.65963138194, 4781.32140186133, 4923.45785956592, 4851.874613326, 
    4797.04288115436, 4877.32098573248, 5200.96937649842, 5446.25232035071, 
    5500, 5343.12737175836, 4751.38004958183, 3649.80765166407, 
    2514.96531355827, 1592.13427519466, 806.119198945454, 429.073855485613, 
    190, 100, 80, 90, 90, 70, -0, -0, -0, -0, -0, -0, 40, 60, 70, 80, 90, 90, 
    -0, -0, 1877.51130615383, 2273.71565894661, 2417.518085942, 
    2672.22454462207, 3152.40875107829, 3517.24190869771, 3827.36991635421, 
    4020.24077474217, 4020.24077474217, 3947.30668182314, 3609.77352896418, 
    3147.8480356343, 2939.90978834303, 2939.90978834303, 3065.78548661781, 
    3132.77515309213, 3375.12421325824, 3580.05415708928, 3738.41374032805, 
    3770.87020520633, 3401.58999935075, 3042.71499317314, 2867.08298528321, 
    2437.4116062552, 2707.76609396034, 2943.14652874087, 3083.47425406967, 
    3073.26640696923, 2974.97128985875, 2901.85858954938, 2857.75401352125, 
    2786.41606762896, 2723.55733096733, 2618.34305728668, 2470.65786246607, 
    2363.73884225747, 2233.26401506668, 2281.00511551577, 2470.85012885614, 
    2758.41088867188, 3288.81683827155, 3603.95711829178, 3897.29707159163, 
    3730.766629041, 4021.58646202477, 4377.66883699158, 4607.68974075311, 
    4987.39500898261, 5202.39869235299, 5319.11204341869, 5233.08646539162, 
    4993.53886326512, 4582.84186018721, 4216.78498758478, 4246.52420182272, 
    4595.8541573611, 4884.15186147549, 5044.3766815079, 5045.03797528777, 
    5024.31988688086, 4985.00952813188, 4961.61881291475, 4914.68603572518, 
    4760.32348776472, 4547.18090028208, 4219.46756567381, 3986.49473290313, 
    3905.78846252809, 3813.52538679381, 3777.20370958049, 3787.19755568141, 
    3878.64645725123, 3953.55006903892, 3949.8403433462, 3822.83937428225, 
    3748.80175078162, 3803.39797042987, 3938.77754269769, 4087.72840545616, 
    4183.76162382327, 4243.83809582861, 4237.41065933828, 4202.2512331351, 
    4115.82976431627, 4036.32232979523, 3993.13225513436, 3964.44559934136, 
    3954.69228998988, 3927.53269438535, 3879.54513101388, 3837.5651079633, 
    3775.96985093827, 3735.49235819346, 3694.09956863997, 3654.681470458, 
    3625.33318610089, 3579.85973403754, 3508.39255117455, 3425.56643795225, 
    3298.89076673688, 3203.12532943881, 3147.54209376608, 3105.00903494538, 
    3112.87900308976, 3162.03188987323, 3248.31508621808, 3366.09020751239, 
    3492.66537051712, 3603.87332563025, 3721.27612304688, 3844.85785310505, 
    3958.52453541711, 4037.09149408501, 4037.09149408501, 4020.79254378777, 
    3939.56395467311, 3869.80718006974, 3791.91777505572, 3748.11273247008, 
    3696.98678626696, 3721.27612304688, 3748.38663413062, 3814.55834295308, 
    3883.45142738743, 3947.54638277622, 4013.14417484927, 4096.45399484948, 
    4184.34740482677, 4284.11484137393, 4419.18185522252, 4560.98528429427, 
    4684.11071776103, 4752.59413281134, 4766.56342419382, 4745.13222089769, 
    4653.15413989085, 4324.58482382753, 3955.70040597996, 3403.0021926752, 
    2466.66776221529, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 2540.0992986978, 3344.89127701425, 3801.14894213316, 
    4195.08036973242, 4425.35841554699, 4527.40374445251, 4650.52120552964, 
    4839.18277979845, 5037.9235120848, 5200.4343094382, 5324.57921044788, 
    5366.86932113542, 5369.52262724763, 5354.30917687506, 5306.26168040122, 
    5243.29277784291, 5143.41858983545, 4989.11708981796, 4798.16967686683, 
    4581.85618050421, 4348.30678812867, 4065.89147763595, 3757.87176526935, 
    3439.3085331511, 3227.00463305649, 3202.68597616808, 3304.21658585486, 
    3466.66988714657, 3641.09005473901, 3770.45695246101, 3868.05442378415, 
    3920.22455177611, 3980.1981127566, 4113.88358570172, 4344.42066312345, 
    4611.86679925756, 4882.15350755015, 5103.79768699509, 5262.59020604933, 
    5431.35431848755, 5500, 5500, 5500, 5476.40614539501, 5381.31666636658, 
    5200.27216788463, 4930.47597621125, 4577.75557347297, 4093.85009922966, 
    3569.05820894546, 3003.10244893368, 2018.27136624409, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 1171.75841196582, 2250, 2250, 2987.744020602, 
    2982.29785149375, 2876.29642943405, 2670.84333571169, 2192.2947123205, 
    -0, -0, 3073.81874474974, 3865.50596760485, 4244.81900129506, 
    4429.20979963361, 4439.95364523435, 4359.24340149026, 4279.96614236261, 
    4107.35588876363, 3676.27877346078, 3119.14304528397, 2403.90820621038, 
    2555.04364325332, 3015.5241601655, 3326.70057069238, 3326.70057069238, 
    3288.6912461234, 3217.50760011534, 3362.65153619088, 3546.76615272805, 
    3775.33970556118, 4013.30022876209, 4329.25564827139, 4665.70398851633, 
    4917.05011168465, 5080.46859034267, 5164.12885961593, 5213.77807425924, 
    5209.74212733364, 5143.41858983545, 5059.66214249196,
  4938.36319448215, 4952.03128819012, 4790.55765486949, 4644.51559719341, 
    4712.94841916801, 4586.62530584034, 4324.27865021182, 4215.46868009883, 
    3501.57949779877, 4643.54707899808, 4780.77618091448, 5256.3666951836, 
    5346.64821734949, 5305.78599375583, 5158.22135649574, 4485.15875541599, 
    4524.52056988161, 4885.01940755142, 5082.18808038991, 5281.55089269713, 
    5355.07185013188, 4873.1619064881, 4753.00792460779, 4783.48534363873, 
    4941.84279595219, 4941.84279595219, 5126.30145342105, 4779.07571895829, 
    4675.33548482761, 4442.010911099, 4767.11289501202, 4669.21682732331, 
    4786.72077626845, 4956.2992162611, 5146.30591395114, 5336.42794316248, 
    5479.96208502713, 5377.24493021528, 4751.38004958183, 3900.32304323373, 
    2593.78786706849, 1857.11162690293, 974.742307018564, 505.043803659173, 
    253.361404418945, 150, 100, 100, 90, 80, -0, -0, -0, -0, -0, -0, -0, 50, 
    70, 80, 90, 90, -0, -0, 1923.41334326407, 2330.55387287496, 
    2705.49464720462, 3255.61393995879, 3335.49707709498, 3540.50877298251, 
    4009.05763982504, 4049.18744100624, 4024.57842026084, 3820.19125279268, 
    3254.31529518305, 2721.17359448501, 2546.3035975955, 2729.74258317126, 
    3159.97449656233, 3169.99662603939, 2951.31545888425, 3479.92890869537, 
    3828.27696481505, 3944.47389131562, 3483.44110383465, 3309.86405150489, 
    2667.94158049595, 2584.65955199799, 2878.25779853487, 3038.80273881526, 
    3038.80273881526, 3009.9432996661, 2877.50994809417, 2849.83515137974, 
    2883.03597704506, 2844.69943735358, 2818.67528656209, 2694.42009833545, 
    2694.42009833545, 2645.26235959542, 2399.98728046216, 2486.33975724372, 
    2885.11465110398, 3031.33276836774, 3362.65764544924, 3500.30693144028, 
    3987.96768699153, 4073.25591099591, 4444.53103472019, 4619.57692354625, 
    4827.49032682229, 5054.99762703953, 5182.36216442919, 5253.03382667717, 
    5161.79680180085, 4906.4036867815, 4041.85917143305, 3532.48138435279, 
    3582.49947945094, 4477.25810145819, 4918.06834314033, 5081.11820449831, 
    5126.05238519283, 5110.18397025516, 5078.40512883347, 5078.40512883347, 
    5053.8018026217, 4927.40744932256, 4697.51455756838, 4403.85510825074, 
    4392.32033320918, 4224.87141153833, 4310.48624346912, 4361.99259735597, 
    4344.85630708721, 4344.85630708721, 4286.45739487234, 4311.93733473737, 
    4152.85954568879, 3993.083186161, 3923.34622082578, 4006.19969118874, 
    4105.23755750869, 4163.52693807315, 4258.07633043667, 4245.34446432785, 
    4223.60228715447, 4095.75190074434, 4010.53519446173, 4009.97713286404, 
    3939.45433923314, 3936.20027379882, 3944.27372106188, 3906.42908019752, 
    3894.65875084573, 3766.36128465078, 3746.01810987184, 3703.66974827996, 
    3663.71094117721, 3644.84413662708, 3614.51160046791, 3579.6136374287, 
    3461.03118879353, 3269.93889890907, 3161.58284719774, 3179.67206522596, 
    3140.35477700321, 3140.12193083941, 3122.33086854763, 3180.78002804977, 
    3317.65484230264, 3460.25421494499, 3590.65328319433, 3708.69954619371, 
    3837.50430224204, 3966.65723543383, 4136.43086312219, 4147.41565957026, 
    4106.01857953561, 4031.1945466833, 3984.82856944387, 3897.96997231054, 
    3826.46812665662, 3768.69399913286, 3697.68400890894, 3732.43476174053, 
    3755.72743432539, 3843.22273696698, 3927.80005675756, 4016.36782560307, 
    4052.66101508359, 4131.11427636261, 4217.48352595958, 4302.54392270554, 
    4456.4288851237, 4597.20875260514, 4740.65269483505, 4740.65269483505, 
    4728.46025511613, 4607.21290571502, 4295.05554282266, 3955.70040597996, 
    2563.39936177336, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 1581.61136303215, 3135.66350385805, 
    3778.76296379547, 4101.6146061721, 4318.52988089467, 4526.86023058006, 
    4615.57111368953, 4933.33590164315, 5153.81989424665, 5358.41359299956, 
    5422.19648100803, 5428.78034372194, 5382.51299992966, 5335.85141819071, 
    5206.59912187907, 5277.23582782817, 5151.22855631407, 5025.67960321167, 
    4812.86508929304, 4603.34361805646, 4352.98117892339, 4137.64043948722, 
    3755.52399784629, 3398.08035893511, 3104.04197761796, 3235.25708336418, 
    3373.58787652753, 3615.87993723466, 3784.54146926086, 3935.29601678296, 
    3959.70372353738, 3974.49563175445, 3866.26308310604, 3845.16982651271, 
    4320.15516109796, 4546.5044581885, 4662.25919283988, 5121.36017958114, 
    5271.50640871299, 5452.24372712278, 5500, 5500, 5500, 5486.40191858117, 
    5399.49790849336, 5223.11988110693, 4958.75989465088, 4616.19577792897, 
    4160.52021729739, 3635.77422304962, 3003.10244893368, 2018.27136624409, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 1171.75841196582, 2250, 2250, 
    2982.29785149375, 2982.29785149375, 2837.93028444651, 3024.41759921419, 
    2487.70974926624, 1544.04810028272, -0, 3242.41021366408, 
    3960.10135754272, 4348.76956723485, 4485.38952592198, 4480.40256147969, 
    4327.46423485733, 4295.16985286639, 4188.98912354307, 3704.06895413281, 
    3324.40509896294, 2450.62181979588, 2487.64161880053, 3015.5241601655, 
    3326.70057069238, 3326.70057069238, 3260.09049179951, 3158.88483692973, 
    3350.16291563405, 3609.74309452673, 3721.27612304688, 3926.55014764471, 
    4280.79807011899, 4648.47693926383, 4898.2078456237, 5088.45391817323, 
    5192.96839517145, 5248.33586134336, 5277.66788917049, 5183.3037318525, 
    5074.46579526224,
  5041.45748418364, 4953.23106523562, 4866.68593981084, 4751.42697163374, 
    4751.42697163374, 4744.23756775728, 4463.67958728863, 4335.33354563713, 
    3983.8227815813, 4535.86022235381, 4858.36721984887, 5214.55136005549, 
    5390.85263362663, 5297.51556636532, 5048.58984881436, 4669.64005415056, 
    4638.84136718881, 4789.46692472072, 5018.2273365821, 5131.03914719227, 
    5111.35457676845, 4850.79968228189, 4766.43317769038, 4859.57302557831, 
    4976.65122011239, 5096.09851119974, 5060.52299361848, 4956.88102326809, 
    4867.60264164018, 4638.77343326813, 4441.61696357712, 4288.27264624545, 
    4394.68579450144, 4640.71264781875, 4857.74648410005, 5143.41858983545, 
    5264.16534063238, 5143.41858983545, 4695.76328563606, 3892.4535442982, 
    2848.80866280136, 2047.13809309956, 1250, 1250, 1250, 240.561416625977, 
    180, 120, 90, 80, -0, -0, -0, -0, -0, -0, -0, 50, 70, 70, 80, 80, -0, 
    770.190877520832, 1923.41334326407, 2330.55387287496, 2683.77380848426, 
    3077.22640044981, 3335.49707709498, 3540.50877298251, 3643.29918040677, 
    3613.53856770945, 3516.15516816456, 3294.61345735061, 3065.78548661781, 
    2721.17359448501, 2640.06400575861, 2692.15704012653, 2904.09554367159, 
    2951.31545888425, 3032.90604852096, 3503.67997515742, 3819.73835535333, 
    3944.65821555356, 3776.11778709742, 3602.68634907351, 2866.33405578437, 
    2609.5182077778, 2849.6412788102, 3038.80273881526, 3054.38397095117, 
    3054.38397095117, 3008.91591987511, 3111.62490203082, 3067.38894505842, 
    3029.22373546945, 2989.97836315402, 2965.1364372857, 2832.6383042203, 
    2685.61127109638, 2476.01839209162, 2593.72315614663, 2780.19843668099, 
    3223.92681861302, 3649.61921404259, 3822.94493103777, 4150.27427017246, 
    4352.47465955445, 4472.0819718012, 4635.30387498498, 4851.55126930362, 
    5028.04038321305, 5099.56519969576, 5031.36469564075, 4919.33769277168, 
    4475.14481996913, 3857.10676880412, 3477.33587176609, 3598.45807866855, 
    4294.17865615644, 4802.95839814511, 5085.28654718102, 5177.99663249337, 
    5190.08513771653, 5176.06028743323, 5183.82894228759, 5082.95120149698, 
    4957.46427089771, 4737.8072900125, 4600.90848752542, 4533.90384444065, 
    4484.28896920877, 4509.49647879075, 4528.55737154832, 4552.59027543899, 
    4551.03417448499, 4564.853048062, 4492.23236919768, 4292.92656753476, 
    4088.02661341309, 3962.19242200561, 3952.77228831498, 4020.49060756897, 
    4103.58166195637, 4194.02506144284, 4198.49942551892, 4176.197139041, 
    4099.52897121509, 4047.41278927426, 4033.70110904626, 4011.50685529843, 
    3995.25414897084, 3959.66136509466, 3917.69359394309, 3886.36630365009, 
    3836.4236200311, 3788.32965267217, 3737.74846186266, 3721.27612304688, 
    3721.27612304688, 3674.09327704433, 3631.02704224907, 3549.75312933356, 
    3423.41676495414, 3342.96327156871, 3289.82359356283, 3230.92735321478, 
    3166.64017585583, 3135.08121840794, 3170.40769326727, 3286.36204913951, 
    3433.79137311609, 3572.22867009597, 3709.44279207017, 3857.96579804337, 
    3995.73377574281, 4142.74920546211, 4178.13913232005, 4151.31699888957, 
    4099.24043345165, 4048.19054086256, 3956.42219706345, 3863.1357219316, 
    3774.08742918745, 3690.05687148416, 3694.99119522707, 3761.78580087913, 
    3851.91649833731, 3943.01965871306, 4027.25796033643, 4082.71703674391, 
    4141.19297800955, 4229.33598808477, 4323.34345987735, 4424.42081680806, 
    4531.7899469825, 4628.98181974321, 4685.76428256175, 4691.87283863985, 
    4461.56603760972, 4130.29982459989, 3525.63102828144, 2373.53437910444, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 2689.00617627103, 3476.52591375365, 3915.68757590321, 
    4208.75516994972, 4492.15744919687, 4643.3040360774, 4932.93457800406, 
    5187.81366770814, 5354.65354984761, 5422.06637090714, 5450.04914717328, 
    5447.12984537784, 5418.21317368935, 5360.45488764167, 5278.16122739706, 
    5166.14894807044, 5021.85831390855, 4841.32507367684, 4637.7326249502, 
    4397.37806189182, 4101.45117547948, 3781.1838499831, 3482.047104524, 
    3240.64022432729, 3247.90056559631, 3373.58787652753, 3598.98690393819, 
    3808.55074527711, 3986.50386689125, 4065.89147763595, 4078.24098130854, 
    4079.0419042854, 4121.20726873034, 4373.61924431739, 4651.55051485441, 
    4805.77975341314, 5074.35665528558, 5261.15675527633, 5440.37262497232, 
    5500, 5500, 5500, 5485.84960528423, 5381.07248951246, 5208.51142993459, 
    4957.59432887365, 4629.20199370764, 4198.27200705086, 3603.88416681283, 
    2981.04638605955, 2177.23583761252, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    1522.00591772311, 2250, 2250, 2835.39492400831, 3017.8268561612, 
    3045.22258240696, 2942.3201308378, 2708.30530998545, 2329.81849342788, 
    2486.26201225781, 3334.23689708705, 3934.03186845636, 4290.83021722284, 
    4474.52272723998, 4438.39975859649, 4302.65398770439, 4213.08431389183, 
    4100.11363174107, 3704.06895413281, 3085.85267961117, 2399.70470884378, 
    2197.50107060228, 2758.41088867188, 3235.58503017594, 3348.67952842066, 
    3348.67952842066, 3286.31681530864, 3411.49659423892, 3581.40240965815, 
    3721.27612304688, 3830.43057282964, 4132.85079232756, 4494.4519865161, 
    4844.53335567439, 5063.08565247005, 5199.8346881226, 5265.01108132914, 
    5296.99109048656, 5239.81645549532, 5156.85654874175,
  5094.2050458072, 4997.76825872152, 4905.77831697895, 4831.05600722653, 
    4751.42697163374, 4744.23756775728, 4656.42282295591, 4513.55275516175, 
    3983.8227815813, 4536.82829508058, 4867.85604164201, 5151.21025814361, 
    5354.15533001993, 5274.77754415436, 5086.78831957652, 4883.16012415236, 
    4700.71822477685, 4761.98136564624, 4978.00301577541, 5007.03588399446, 
    4981.97837897542, 4904.49199053912, 4900.72488077343, 4865.7852708563, 
    4810.78245774324, 4991.39642932177, 5091.8085512988, 4987.30028079769, 
    4877.33273649559, 4590.95199768278, 4355.16057107273, 4200.88925768443, 
    4178.1898568776, 4383.50767635943, 4573.57776514517, 4876.27203528544, 
    4974.39820296112, 4832.20157562459, 4419.18185522252, 3721.27612304688, 
    2807.06764207379, 2063.27720478932, 1250, 1250, 1250, 1250, 180, 120, 90, 
    80, -0, 40, 40, 50, 50, 50, 50, 50, 60, 70, 70, 70, -0, 770.190877520832, 
    1562.92689347154, 1980.39634693846, 2443.73153365325, 2828.36174375482, 
    2959.16806881348, 3001.21382332797, 2979.26968770345, 2887.06093194787, 
    2744.96863938093, 2573.91974904123, 2656.8181650283, 2656.8181650283, 
    2732.29259756555, 2729.02831349596, 2894.51610295153, 2870.61648374515, 
    2986.19632109408, 3543.70255366377, 3867.16960604271, 3947.83339327582, 
    3792.47290416295, 3587.55642736927, 2777.40983211065, 2759.72893521272, 
    2923.13806519825, 3038.80273881526, 3054.38397095117, 3054.38397095117, 
    3008.91591987511, 3330.73335219819, 3322.933615373, 3192.29622692419, 
    3323.46027760103, 3268.85303378237, 2988.61624316413, 2685.61127109638, 
    2740.96469323867, 2889.73508724633, 3232.82895584059, 3560.73689372535, 
    3876.78683917395, 4086.05019788389, 4230.61584402675, 4353.26829547624, 
    4483.73973357784, 4679.8436899619, 4885.81426305237, 4973.10921484458, 
    4978.25418032183, 4876.3950080527, 4564.44204536764, 4109.22139299235, 
    3664.06786445573, 3349.88191882324, 3526.0676337227, 4198.71607468009, 
    4779.75252921983, 5071.65470009082, 5213.16523394079, 5264.14027432547, 
    5283.63129929734, 5246.00750842457, 5123.87277886758, 4975.32498289319, 
    4742.01127806868, 4686.2535624883, 4650.70761562767, 4657.22793319948, 
    4713.63008654024, 4728.55090559784, 4718.03459567224, 4705.95439096313, 
    4662.1951853395, 4565.10136343707, 4365.04893234209, 4084.23527418666, 
    3918.16631085422, 3864.5596883224, 3920.55270680981, 4045.79400518843, 
    4152.78301277781, 4179.81238826119, 4166.30097065688, 4118.61003560137, 
    4047.41278927426, 4052.73783003426, 4052.73783003426, 4034.07833166995, 
    3978.3457180407, 3934.96136710821, 3885.81486618723, 3854.50793282605, 
    3797.33966515674, 3770.980830846, 3774.38274183304, 3791.35733216571, 
    3791.43246688081, 3747.96688290889, 3678.42939166811, 3587.86350087068, 
    3490.63858749391, 3403.30668393832, 3320.3547135238, 3221.67018748551, 
    3154.19155938571, 3153.7138221073, 3252.68109701337, 3406.22887490465, 
    3551.81937193178, 3693.89977647834, 3861.34377780062, 4010.85259667751, 
    4156.91972992379, 4205.33351788443, 4192.26655841114, 4158.75513885827, 
    4105.31489953476, 4003.66293889756, 3909.12977562016, 3793.50883695786, 
    3708.7765377494, 3697.79313862188, 3772.74335044611, 3863.80730132704, 
    3958.14007017829, 4049.69455795193, 4111.0067036295, 4170.09192125605, 
    4243.74460410173, 4324.08334790045, 4407.87633911928, 4492.83017957339, 
    4565.60822190238, 4626.30422628209, 4602.48554104308, 4294.87899090084, 
    3918.13716506946, 2936.265125934, 2009.32352529971, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    3101.78388261717, 3690.17856410796, 4065.89147763595, 4452.06765221688, 
    4686.80184362656, 5005.21798541142, 5219.43581625254, 5362.61895385608, 
    5439.69596737638, 5466.0989693728, 5474.37726961716, 5452.14637406153, 
    5417.75361996753, 5316.33724265876, 5193.69511929956, 5027.70235930194, 
    4845.43961709801, 4628.52485147203, 4396.85302742195, 4127.2189076176, 
    3795.58418271572, 3497.23941274529, 3260.82107729789, 3199.29865562509, 
    3331.22965121022, 3556.47175633318, 3817.57801322842, 4002.30762516286, 
    4113.21524020134, 4127.81623418371, 4162.09937227772, 4238.85706321548, 
    4434.51337349289, 4693.41119588839, 4854.35596670509, 5001.0377570304, 
    5220.21654751018, 5446.14158949426, 5500, 5500, 5500, 5483.42736164662, 
    5365.64160566526, 5190.05182548343, 4949.01807185483, 4649.8365706384, 
    4214.55062790976, 3610.72405274501, 2958.08020056065, 2177.23583761252, 
    0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 1575.89572955051, 2250, 2250, 
    2801.79600567705, 3164.45825204639, 3263.22434985506, 3254.59696626337, 
    3101.70854465349, 2959.26170951102, 2895.83216901697, 3334.23689708705, 
    3894.71291581909, 4269.03467701147, 4372.95994161556, 4372.95994161556, 
    4233.72541127596, 4133.35731103926, 3980.73892599243, 3550.29193196041, 
    2853.39625272245, 2191.85384798669, 1841.6107979499, 2413.34888528194, 
    3091.55979337995, 3420.19428843832, 3431.63611545133, 3286.31681530864, 
    3453.7463327077, 3559.70614606956, 3644.01237958072, 3658.75881226187, 
    3939.84239410192, 4364.0498511475, 4779.07571895829, 5046.73379237748, 
    5210.13285962137, 5303.05290022056, 5321.61708810168, 5275.42579470477, 
    5201.24163169666,
  5131.3, 5032.2, 4949.5, 4903.4, 4837.8, 4850.5, 4736.6, 4598.5, 3954.4, 
    4589.9, 4892.4, 5143.41845703125, 5297.1, 5274.5, 5129.9, 4953.2, 4847, 
    4882.1, 5028, 5020.3, 5053.6, 5048.8, 5029.8, 5009.9, 4892.4, 4880, 
    5037.8, 4923.7, 4698.3, 4419.181640625, 4355.16057107273, 
    4200.88925768443, 4178.1898568776, 4383.50767635943, 4573.57776514517, 
    4573.57776514517, 4065.89147763595, 4439.94375794645, 4608.57571467985, 
    3721.27612304688, 1890, 980, 685.391009172411, 1250, 1250, 1250, 1250, 
    110, 90, 80, 80, 70, 40, 50, 60, 60, 50, 50, 60, 60, 50, 40, -0, 190, 
    1406.18801489997, 1381.84224278682, 1666.74311165122, 2196.32692357124, 
    2196.32692357124, 2022.9883441464, 1182.87476765165, 600.077251875481, 
    425.785466617812, 2246.6, 2310.8, 2345, 2403.1, 2674.7, 2723.2, 2723.2, 
    2820, 3098.8, 3564.9, 3700.9, 3633.9, 3332.8, 2825.3, 2860.7, 3121.3, 
    3336.7, 3485.3, 3560.1, 3579.5, 3819.4, 3832.1, 3756.2, 3827.1, 3727.8, 
    3494.1, 3151.2, 3179.3, 3387.2978515625, 3661.1, 3860, 4036.6, 4164.2, 
    4245.3, 4319.3, 4451.5, 4644.5, 4784.4, 4779.07568359375, 4701.7, 4572.9, 
    4350.6, 3970.7, 3567.3, 3330.9, 3558.6, 4210.4, 4785.6, 5092.5, 5241.6, 
    5278.4, 5500, 5225.1, 5107.5, 4893.7, 4760.5, 4697.5, 4669.5, 4728.5, 
    4779.07568359375, 4790.8, 4779.07568359375, 4757.1, 4687.6, 4538.6, 
    4365.04893234209, 3995.8, 3792, 3700.9, 3892, 4045.7, 4165.3, 4212.2, 
    4204.4, 4183.6, 4145.6, 4144.1, 4137.2, 4107, 4038.9, 3988.6, 3939.6, 
    3901.9, 3859.7, 3846.4, 3867.4, 3891.6, 3917, 3893.7, 3830.2, 3735.9, 
    3632.9, 3518.2, 3398.5, 3288.1, 3192.7, 3159.5, 3229.8, 3368, 3514.4, 
    3655, 3829.3, 3982.5, 4147.6, 4219.1, 4230.1, 4187.6, 4131.6, 4034.8, 
    3927.7, 3810, 3727.8, 3693.4, 3791.3, 3897.1, 3990.6, 4079.7, 4137.9, 
    4195.3, 4259.4, 4325.5, 4393.9, 4468.2, 4531.4, 4579.8, 4450.9, 4112.7, 
    3493.4, 2280.3, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 1346.80157430838, 3389.8, 3946.7, 
    4393.3, 4713.1, 5036.7, 5221.9, 5354, 5435.4, 5483, 5487.2, 5476.1, 
    5447.5, 5353.5, 5235.4, 5050.6, 4859, 4634.6, 4393.5, 4111.9, 3800, 
    3483.4, 3226.9, 3105.7, 3186.1, 3462.1, 3742.5, 3957.8, 4350.01084157075, 
    4161.3, 4208.5, 4292.9, 4476.1, 4679.6, 4846.8, 4986.2, 5133, 5500, 5500, 
    5500, 5500, 5500, 5333.5, 5156.4, 4928.1, 4637.9, 4209.3, 3566.6, 2817.5, 
    2045.9, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 1050, 2250, 2250, 3032.5, 
    3450.40774825414, 3547.14762441652, 3617.38898014786, 3617.38898014786, 
    3586.89855590781, 3619.52106871343, 2897.853093021, 3817.8, 4178.7, 
    4309.6, 4271.1, 4123.9, 3919.9, 3784.2, 3321.8, 2611.4, 1117.9, 729.7, 
    2316.1, 3068.9, 3457.9, 3507.1, 3366.9, 3472.5, 3542.6, 3559.7, 3407.6, 
    3726.1, 4193.3, 4691, 5006.6, 5198.2, 5299.4, 5333.1, 5301.3, 5230.9,
  5168.4041537152, 5066.5966470579, 4993.23978968884, 4975.76044694226, 
    4924.19850429116, 4956.66946273908, 4816.86945301888, 4683.36399530974, 
    3925, 4642.90350774659, 4916.9752248878, 5119.25200792029, 
    5240.12385551799, 5274.28014773672, 5172.93958055771, 5023.24664144141, 
    4993.31819529193, 5002.28980373868, 5078.06489915659, 5033.58020828136, 
    5125.25073104055, 5193.03919824137, 5158.91331096019, 5154.00075313556, 
    4974.01803373829, 4768.53188595288, 4983.83156231898, 4860.13242563934, 
    4519.18559984027, 4231.11477874334, 3946.97306662225, 3721.27612304688, 
    3555.50551888782, 3489.07465246811, 3556.37130658771, 3787.24922036347, 
    3818.1229098173, 3662.29800943104, 3294.45618235304, 2721.77518107038, 
    1890, 1890, 1890, 0, 1250, 1250, 1250, 1250, 447.69390685827, 
    370.154968261719, 270.610395222517, 190, 130, 90, 70, 60, 60, 50, 50, 50, 
    50, 50, 0, 190, 962.24776583742, 1373.06821198615, 1666.74311165122, 
    2033.39408104555, 1967.48950326866, 1732.49850931692, -0, 
    1746.58497734966, 2097.58841179977, 2519.30373549249, 2764.81843798564, 
    2833.1001030491, 2873.81565733392, 2620.42525091447, 2607.04401189127, 
    2575.80557871653, 2653.80337120715, 2653.80337120715, 3262.64426151785, 
    3453.99680722876, 3475.31776723964, 3078.01260881568, 2873.11425317972, 
    2961.68495409187, 3319.4592264436, 3634.52626150024, 3916.14507775483, 
    4065.89147763595, 4150.15117368846, 4308.05080097564, 4341.27593774945, 
    4320.15522485821, 4330.7766090106, 4186.73998903889, 3999.50723772002, 
    3616.84680258864, 3617.6619180194, 3880.52560687722, 4089.40634881211, 
    4159.30314550682, 4196.46493377798, 4242.40044959366, 4260.02459885591, 
    4285.36124689015, 4419.18185522252, 4609.12542442931, 4683.06147463124, 
    4567.2989167888, 4425.11309499512, 4269.43569997926, 4136.69069026453, 
    3832.23660622585, 3470.47681732335, 3311.82071392678, 3591.04678324455, 
    4222.15820641331, 4791.50315309507, 5113.44272799958, 5269.93877256461, 
    5292.61231769255, 5317.31607108133, 5204.11234526658, 5091.20851193389, 
    4812.12151257607, 4779.07571895829, 4708.72441781839, 4688.19359613195, 
    4799.85384817479, 4832.54625895363, 4852.97600677043, 4839.82685348893, 
    4808.27309614982, 4713.03031765455, 4512.18688694958, 4193.71774852098, 
    3907.45420427209, 3665.92296450681, 3537.30458794967, 3863.48279489608, 
    4045.58139590202, 4177.84656092431, 4244.66483550655, 4242.42154765261, 
    4248.66228666475, 4243.76789940926, 4235.55857978146, 4221.60351658737, 
    4179.92332443252, 4099.4246291591, 4042.16133242119, 3993.29653795138, 
    3949.20084399853, 3922.0686687991, 3921.89230608033, 3960.3588550541, 
    3991.90161029925, 4042.5877490038, 4039.52194151897, 3981.96488127011, 
    3883.85307105669, 3775.245445821, 3633.18552872974, 3476.57006203845, 
    3354.53963381203, 3231.22760486652, 3165.25388450374, 3206.9869702095, 
    3329.74730089257, 3476.98832426168, 3616.12479881334, 3797.2040219255, 
    3954.20374562253, 4138.27265985072, 4232.92527179893, 4267.9381515331, 
    4216.51420132043, 4157.87974887032, 4044.08928875994, 3946.26910997416, 
    3826.46735152407, 3746.85083818481, 3688.9730499142, 3809.8888969488, 
    3930.32916018171, 4023.05828299163, 4109.7869914027, 4164.85507722184, 
    4220.51019859977, 4275.05542219352, 4326.90772980739, 4379.89429874486, 
    4443.6641246688, 4497.2652648513, 4533.38228900712, 4299.41242418858, 
    3930.43824311445, 3068.72451800475, 1624.42864963155, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    0, 3089.4885168817, 3827.51375394589, 4334.60996247262, 4739.45501861666, 
    5068.09649084134, 5224.45089363377, 5345.43892941164, 5431.11366276773, 
    5500, 5500, 5500, 5477.33846254847, 5390.60733429202, 5277.0561847089, 
    5073.53713069016, 4872.64676637801, 4640.69987649039, 4390.12461781063, 
    4096.51539403799, 3804.48659025377, 3469.48753765754, 3193.00559675806, 
    3012.11517214948, 3041.0011064085, 3367.76370419449, 3667.45746231496, 
    3913.35503036803, 4092.79334715687, 4194.87204842616, 4254.83924244087, 
    4347.03602772875, 4517.71482362791, 4665.7599151078, 4839.20536113254, 
    4971.39103081866, 5045.71089082394, 5369.23214240698, 5500, 5500, 5500, 
    5445.87386175295, 5301.45552151846, 5122.70488309205, 4907.16834681443, 
    4625.86927408133, 4204.11053592294, 3522.50510385056, 2676.8384704844, 
    1914.49516980276, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 1799.28378123357, 
    2250, 2250, 3263.21148289574, 3457.67348409005, 3562.29945368972, 
    3633.69231602058, 3617.38898014786, 3586.89855590781, 3544.10988090116, 
    3332.52182629931, 3740.97181724108, 4088.38782540114, 4246.28444045303, 
    4169.23322162298, 4014.15425440938, 3706.4716807934, 3587.75635165566, 
    3093.34395690737, 2369.42495846932, 1643.98141881264, 1617.88810259288, 
    2218.79526570893, 3046.24805213255, 3495.59056603977, 3582.48421664866, 
    3447.45345738227, 3491.34664937496, 3525.4567366724, 3475.44213172107, 
    3156.43621874857, 3512.28496062241, 4022.48413622147, 4602.82571040104, 
    4966.50871409275, 5186.2477569751, 5295.6733081685, 5344.50301797447, 
    5327.17952300628, 5260.63336715414,
  5187.90451235258, 5055.72446684596, 5012.06839280879, 4977.55114314676, 
    4943.98517371624, 5004.69399766336, 4858.43157596325, 4719.97528718838, 
    3926.02196501208, 4637.58945939762, 4916.50089649773, 5119.25200792029, 
    5240.10449921716, 5219.6675925073, 5210.5739424129, 5075.82323203556, 
    5122.06456163685, 5079.51811445742, 5156.2251054844, 5216.0378153096, 
    5236.74861357633, 5307.81203219523, 5304.07527987095, 5204.31497503596, 
    4988.17295949033, 4766.58869204818, 4751.86865772491, 4440.72814060327, 
    3970.99394338184, 3556.73335939334, 3192.48287306945, 3133.16880026756, 
    2988.89513613811, 2925.92611968449, 3090.58946816395, 3161.06723765257, 
    3109.71391650843, 2889.05767922219, 2529.81289303451, 1890, 1890, 1890, 
    2085, 2085, -0, 1250, 1250, 1250, 803.91847147382, 672.809708258495, 
    505.281363965325, 240.561416625977, 190, 110, 80, 60, 60, 50, 50, 50, 50, 
    50, 0, 190, 683.282409667969, 1185.46767400173, 1185.46767400173, -0, -0, 
    0, 425.785466617812, 1861.85711054023, 2083.38470330905, 
    2486.32563819725, 2913.29209524067, 2937.33151363858, 2865.46124004852, 
    2722.7129789794, 2503.87762478546, 2233.69370246163, 2159.95161813917, 
    2414.44693350829, 3189.61663642711, 3363.16895996019, 3363.16895996019, 
    3186.26163638822, 3121.58545426414, 3257.33774527363, 3591.04060314314, 
    3912.76979780307, 4182.0154376088, 4444.03949508165, 4635.57892449908, 
    4719.02721495743, 4729.69320112879, 4705.12128944456, 4615.43721283197, 
    4446.72104901239, 4297.1759356774, 4085.52459805358, 4142.92079269027, 
    4333.42107781393, 4524.88661764304, 4598.83655913123, 4545.52366967626, 
    4397.16005130937, 4324.44931928886, 4271.13372729575, 4265.37153301421, 
    4481.61500507756, 4599.45988716781, 4475.85647427606, 4304.16133445129, 
    4096.07041285614, 3908.30940566935, 3788.98319945077, 3509.78592367029, 
    3311.82071392678, 3795.51328887442, 4274.01295839493, 4834.00083691422, 
    5126.66649638236, 5239.50875081638, 5296.1361431906, 5289.63264453565, 
    5224.77631714143, 5025.63907356059, 4804.13047659461, 4779.07571895829, 
    4692.82875848606, 4794.76060198641, 4846.42823407842, 4892.88710573532, 
    4906.5152297123, 4896.50918082585, 4825.40812263923, 4674.37480645706, 
    4419.18185522252, 4101.92368456849, 3737.18428089039, 3502.06471475586, 
    3599.70401141708, 3932.88022109365, 4129.56395641192, 4283.0407996989, 
    4361.03515125196, 4384.89256969429, 4387.00528549404, 4377.12386057122, 
    4366.07423194883, 4353.97005165412, 4294.43384641767, 4213.81752163564, 
    4138.31738252081, 4076.40172477886, 4043.18318015056, 4021.73396093868, 
    4017.13598101548, 4069.57387323551, 4114.7108363936, 4158.16880260351, 
    4161.27372171545, 4110.68419748784, 3999.66360706191, 3890.62218854052, 
    3737.209621095, 3563.34079393574, 3424.33079475609, 3286.32825295191, 
    3195.80842668763, 3204.3497675451, 3296.33966407863, 3431.20061010587, 
    3554.44932973563, 3724.2883762643, 3891.61040906858, 4090.16763053796, 
    4214.94666179072, 4232.96750215356, 4219.60392430185, 4155.16053605236, 
    4044.08928875994, 3940.11153230088, 3840.28874290029, 3779.69261522085, 
    3776.79110500813, 3863.37332626392, 3986.55876159393, 4041.45872803633, 
    4114.76312005679, 4170.15038677124, 4224.68460619212, 4269.9329403566, 
    4326.07438534647, 4378.1085225511, 4419.18185522252, 4462.81321237507, 
    4420.36230863986, 4130.77973427334, 3661.07646587327, 2397.99992824023, 
    1624.42864963155, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 2555.02503647793, 
    3557.97695993746, 4257.89221382984, 4710.89924494458, 5046.83222588913, 
    5237.38286775488, 5333.63170331469, 5434.6036596576, 5500, 5500, 5500, 
    5500, 5431.78838413653, 5292.52157452565, 5062.04331648435, 
    4812.668365175, 4580.59109511862, 4349.92773882039, 4078.20988315531, 
    3788.23948374484, 3469.16159014493, 3183.79840620809, 2973.66210912785, 
    3041.0011064085, 3305.81293865055, 3588.13817528936, 3799.74607693014, 
    4000.29829388452, 4177.53409546605, 4286.92376962579, 4376.96136807494, 
    4505.14957081758, 4594.02529106301, 4765.26321243419, 4903.67360472501, 
    5045.71089082394, 5279.32984162847, 5495.76723854536, 5500, 5500, 
    5402.74235847846, 5246.34355677494, 5053.4191933554, 4841.30765204428, 
    4562.91293532221, 4147.59021914647, 3431.72647291609, 2565.65644664787, 
    1768.00643635456, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 2127.37502497806, 
    2592.10906889378, 3039.89768335552, 3458.51917848896, 3634.92347883241, 
    3641.51851110525, 3641.51851110525, 3735.76825295397, 3797.01341147303, 
    3760.98766295069, 3332.52182629931, 3641.92048689487, 4050, 4050, 
    4014.50997436057, 3860.23388291303, 3597.93888450641, 3374.14146243877, 
    2833.63091782338, 2149.94877114536, 1643.98141881264, 1906.02833745084, 
    2453.20496801585, 3184.23848284421, 3584.09954569159, 3662.49595156207, 
    3555.64542220448, 3512.47711493958, 3490.18809490393, 3369.36770812735, 
    3156.43621874857, 3246.82303122399, 3733.71169713187, 4456.3757128343, 
    4909.33345747891, 5170.15628834386, 5291.00956338184, 5338.70265122471, 
    5335.89537646666, 5276.39382174384,
  5181.1, 5074.6, 5021.7, 4989.4, 4954, 5024.9, 4908.4, 4756.6, 4217, 4595.7, 
    4890.8, 5071, 5206, 5198.9, 5177, 5116.4, 5116.4, 5113.5, 5183.2, 5500, 
    5500, 5289.3, 5207.9, 5023.7, 4758.7, 4766.58869204818, 4204.41465191137, 
    2675.28681027879, 3094.16637163852, 3226.48378690357, 2157.24306327261, 
    2008.72559722242, 1637.32729792239, 1846.62237651059, 1846.62237651059, 
    1292.80751861564, 913.921661605496, 335.502712964576, 335.502712964576, 
    -0, 629.751742867894, 1890, 2085, 2085, 0, -0, 1250, 1844.48734148472, 
    1844.48734148472, 1520.25594230878, 816.056051104196, 240.561416625977, 
    240.561416625977, 150, 90, 60, 60, 50, 50, 50, 40, -0, -0, 40, 130, 
    534.285534499501, 534.285534499501, -0, -0, 425.785466617812, 930.5, 
    1383.3, 1451.8, 2453.3, 3019.7, 2956.4, 2690.8, 2320.8, 2191.85375976562, 
    1981.1, 2036, 2351.2, 2933.6, 3236.8, 3349.7, 3341.3, 3374.7, 3465.4, 
    3736.8, 4072, 4397, 4669.6, 4859.1, 4942.4, 4941.7, 4897.4, 
    4779.07568359375, 4604.9, 4440.6, 4355.9, 4490.1, 4690.9, 4861.2, 4911.8, 
    4833.9, 4655.7, 4531.9, 4371.9, 4423.4, 4579.2, 4640.8, 4538, 4340.7, 
    4116, 3906.5, 3828.4, 3632.8, 3559.9, 3936.2, 4364.1, 4890.8, 5153.1, 
    5243.8, 5295.9, 5260.4, 5164.9, 5001.1, 4838.6, 4784.9, 4779.07568359375, 
    4871.8, 4923.2, 4971.7, 4954.7, 4898.4, 4785.9, 4610.6, 4349.1, 4027.8, 
    3640.8, 3565.5, 3735.5, 4014.8, 4227.5, 4365.4, 4439.9, 4471.4, 4487.2, 
    4480.4, 4467, 4451.8, 4394.4, 4328.6, 4263.2, 4207.3, 4174.9, 4156.7, 
    4140.3, 4176.3, 4200.3, 4223.2, 4221.3, 4176.1, 4082.5, 3972.7, 3823.8, 
    3643.3, 3502.2, 3365.4, 3266.2, 3241, 3277, 3371.9, 3493.5, 3658.5, 
    3826.2, 4002.4, 4140.4, 4157.2, 4155.8, 4102.7, 4010, 3921.5, 3839.2, 
    3800.6, 3825.2, 3903.8, 4003.3, 4065.89135742188, 4117, 4156.2, 4202.4, 
    4234.5, 4289.2, 4332.4, 4369.4, 4369.4, 4272.7, 3975.3, 3210.7, 1355.6, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 3273.7, 4145.8, 4665.3, 5026.8, 5248.4, 
    5354.8, 5500, 5500, 5500, 5500, 5500, 5447.4, 5305.7, 5058.2, 4821.3, 
    4565.4, 4321.1, 4065.89135742188, 3791.5, 3504.1, 3211.7, 3011.5, 
    3065.78540039062, 3277.1, 3552.6, 3747.8, 3990.7, 4184.2, 4331.6, 4425, 
    4509.6, 4570.9, 4668.3, 4779.07568359375, 4918.8, 5500, 5500, 5500, 5500, 
    5348.2, 5177.6, 4976.4, 4749.8, 4453.3, 4016.7, 3282.5, 2466.66772460938, 
    1571.6, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 314.617511966701, 2149.5, 2692.9, 
    3360.25737446712, 3768.93622810457, 3983.95459459646, 3921.05136661691, 
    3847.41453856124, 3999.28525126085, 4003.2375282488, 4003.2375282488, 
    3642.2, 3757.4, 4050, 4050, 3893.7, 3696.5, 3388.2, 3160.8, 2710.4, 
    2207.9, 2015.8, 2310.7, 2789.7, 3387.2978515625, 3673.9, 3673.9, 3593.6, 
    3493.7, 3461.5, 3287.3, 2948.8, 2988.4, 3475.9, 4272.7, 4819.1, 
    5143.41845703125, 5274.5, 5326.1, 5323.9, 5265.5,
  5174.2820040324, 5093.53448274079, 5031.32412711369, 5001.24289593619, 
    4964.01545694401, 5045.15380502534, 4958.39022989562, 4793.27871667127, 
    4507.98737354995, 4553.85444423204, 4865.00741062468, 5022.69480490463, 
    5171.97520431179, 5178.10947185657, 5143.41858983545, 5156.95423727472, 
    5181.0446580032, 5147.56740315732, 5210.17522887161, 5313.75533602431, 
    5358.61058513068, 5270.76321437053, 5111.64881091774, 4843.07818632963, 
    4529.23107612882, 4018.78877115578, 3397.45620067719, 2675.28681027879, 
    2680.60286672558, 2211.46926623023, 1839.23639879832, 1639.94355960321, 
    1460.29140266812, 1413.7336373015, 40, 40, -0, -0, -0, -0, -0, 0, 2085, 
    2085, 2134.8402921202, 2098.19323649997, 1913.88638739938, 
    1915.4062612279, 1844.48734148472, 1616.86360533153, 1239.4930620529, 
    240.561416625977, 253.361404418945, 253.361404418945, 170, 80, 60, 50, 
    40, 40, 40, -0, -0, 40, 130, 130, -0, -0, 1791.02786294536, 
    2071.500807947, 2251.26159755485, 2704.79311682456, 3220.29267164657, 
    3220.29267164657, 3126.12454940494, 2975.48456357001, 2516.16770520344, 
    1918.82941677571, 1870.47968516987, 1728.48145863056, 1912.136932983, 
    2287.9206460295, 2677.56521469092, 3110.40648977891, 3336.27003062899, 
    3496.2825074199, 3627.8183883731, 3673.50901150173, 3882.64846354988, 
    4231.1804777743, 4611.94662563674, 4895.23049951531, 5082.68358677615, 
    5165.67334873984, 5153.65505910849, 5089.65746631882, 4939.74334043244, 
    4763.04815321214, 4584.04091141102, 4626.3039792622, 4837.31685584943, 
    5048.28828277932, 5197.42661431676, 5224.77917225443, 5122.37067896477, 
    4914.27143248412, 4739.30234747056, 4472.72120468171, 4581.48517472839, 
    4676.85726654754, 4682.11413480593, 4600.17948311141, 4377.22180230683, 
    4135.84911480692, 3904.77384022276, 3867.8450151695, 3755.74527207632, 
    3808.03451729594, 4076.95239907567, 4454.09755069115, 4947.50829092729, 
    5179.59022664199, 5248.02098210376, 5295.59425058188, 5231.14701820231, 
    5105.05252911644, 4976.56636651047, 4873.09095531574, 4790.69680931402, 
    4860.47512201248, 4948.74451714821, 4999.97234033085, 5050.56399728766, 
    5002.90730182579, 4900.30958473678, 4746.40976876996, 4546.89459978581, 
    4279.07492318667, 3953.61441918428, 3544.39161378756, 3628.88218037055, 
    3871.37873466789, 4096.64272545584, 4325.45575109581, 4447.67988636596, 
    4518.76896874635, 4557.83545569619, 4587.49274217876, 4583.70312528793, 
    4567.93910050369, 4549.69159276972, 4494.3186551172, 4443.32474889653, 
    4388.0334131191, 4338.13047570784, 4306.63174851729, 4291.58087545501, 
    4263.55793009286, 4282.92672975838, 4285.83167813716, 4288.28183515107, 
    4281.23692034336, 4241.46326248961, 4165.28543025466, 4054.8187456606, 
    3910.34506036945, 3723.21355549492, 3580.03650994424, 3444.47313364249, 
    3336.51867620416, 3277.56662665306, 3257.61763061084, 3312.53329064718, 
    3432.55096943619, 3592.70011219997, 3760.87290388113, 3914.54219244254, 
    4065.89147763595, 4081.52673288328, 4091.89731523047, 4050.19641652829, 
    3975.82040569307, 3902.9223550996, 3838.05188181024, 3821.56606301982, 
    3873.7068842486, 3944.21029942124, 4019.9945594478, 4074.29526397829, 
    4119.21925728133, 4142.2247357176, 4180.09691555319, 4199.11838506285, 
    4252.33345767977, 4286.77778089245, 4319.53643112866, 4363.79177768095, 
    4124.98040765195, 3819.76259632568, 2760.31132761371, 313.25901422206, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 2989.46597392062, 4033.69336387265, 
    4619.7973363789, 5006.6811290045, 5259.34996520822, 5375.93869409147, 
    5478.77966453167, 5500, 5500, 5500, 5500, 5462.92170268333, 
    5318.9369582857, 5054.39682117382, 4829.88949626886, 4550.23302631214, 
    4292.25370634688, 4047.63049549761, 3794.73738266705, 3539.10586310883, 
    3239.65138315649, 3049.39129002759, 3074.70664515527, 3248.41220043725, 
    3517.02682453804, 3695.85907237597, 3981.10623388679, 4190.77294543225, 
    4376.20374824368, 4473.0795000122, 4514.0489833121, 4547.7762576593, 
    4571.40076372944, 4649.89298683843, 4791.92811291014, 5032.06562726864, 
    5272.4588125479, 5416.68753811226, 5405.72967828517, 5293.59197380116, 
    5108.88842082044, 4899.31688917097, 4658.3654198042, 4343.6838109716, 
    3885.80844441777, 3133.34304862038, 2358.7079556184, 1375.28154311486, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 1369.95677481273, 2171.54833350865, 
    2793.72835699147, 3360.25737446712, 3749.65584403881, 3921.05136661691, 
    3979.56587404503, 3871.62213703227, 3911.64844771242, 4003.2375282488, 
    4003.2375282488, 3951.93150991955, 3872.86986360505, 4050, 4050, 
    3772.9068996789, 3532.80864248176, 3178.48297195721, 2947.39783651585, 
    2587.08487952067, 2265.90841315553, 2387.64490855176, 2715.29940938716, 
    3126.22311702996, 3571.35177009526, 3763.73319094506, 3765.52185718669, 
    3631.52138769039, 3474.95838995603, 3432.74021896918, 3205.13762783879, 
    2741.18857482865, 2729.88525400195, 3218.09365520776, 4089.04704242326, 
    4728.88469105383, 5106.42252904773, 5257.92855732028, 5313.43353519664, 
    5311.95101632689, 5254.55724631176,
  5173.74598346608, 5099.6905916615, 5027.76517549649, 4993.27565356694, 
    4954.06914001258, 5038.63976751539, 4967.88797102306, 4797.83867776249, 
    4537.00042410577, 3925, 4779.07571895829, 4958.57346077224, 
    5095.22827619, 5125.18446393655, 5130.8453524079, 5143.41858983545, 
    5143.41858983545, 5144.47670656859, 5188.2435392659, 5283.60162369075, 
    5257.56966711566, 5024.99097803421, 4779.07571895829, 4350.82979716766, 
    3864.85980216922, 3178.32996124153, 2551.73793897515, -0, -0, -0, -0, -0, 
    -0, -0, 260, 260, 543.62711826946, 718.579702303184, 900.06081491837, 
    1590.94665536754, 1590.94665536754, 1867.56750111359, 2149.3838640566, 
    2428.32567191327, 2652.97025037021, 2652.97025037021, 2556.6584731516, 
    2535.5110626211, 2488.93341400133, 2311.56181338202, 1855.93698466145, 
    -0, 425.785466617812, 425.785466617812, 230, 130, 60, 50, 0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 1684.35603970423, 2423.67666505251, 2942.40047209745, 
    3110.89223808053, 3525.83363354396, 3694.52495345339, 3694.52495345339, 
    3434.09515031485, 2816.9391518884, 2178.45215143225, 1782.77547438591, 
    1738.75447196002, 1808.306182718, 2054.94248553819, 2287.9206460295, 
    2657.70459665775, 3162.61714890441, 3387.2978515625, 3447.64097262201, 
    3555.24804859467, 3697.44924290024, 3916.57240363106, 4237.97280151317, 
    4598.1720284281, 4887.64971863954, 5129.30569049142, 5237.62207919427, 
    5240.93933133432, 5164.57165686985, 4960.43786683703, 4807.81894633368, 
    4623.74306069605, 4816.14027871506, 5006.88537774874, 5226.3520678127, 
    5396.53082904814, 5416.68265814875, 5325.26493407107, 5165.54355627733, 
    4971.53930429083, 4832.28538236691, 4804.07080838031, 4828.58286618232, 
    4893.20821686681, 4805.99260922264, 4492.04781412932, 4216.12955284054, 
    3970.58836123146, 3932.11648671612, 3905.30764182302, 4027.06983309652, 
    4276.8216644608, 4582.56035225767, 4978.79378835645, 5205.01447401956, 
    5268.99216492584, 5227.2529108236, 5180.46915780931, 5074.93265731879, 
    4969.18688438806, 4881.65882405234, 4800.97966818745, 4939.76095033281, 
    5005.67996472797, 5052.75874281431, 5048.99420274501, 4955.8144872168, 
    4843.06133668679, 4689.24401234459, 4507.25495225582, 4285.99370527588, 
    3996.6669209336, 3686.73408456288, 3796.72870975241, 3983.19726383759, 
    4212.89152273508, 4394.62876832401, 4484.34300004978, 4571.51902558505, 
    4607.23879958672, 4634.87242550214, 4630.80093172701, 4610.73860900782, 
    4580.45173722244, 4538.80718154908, 4499.73362496728, 4438.0566905371, 
    4419.18185522252, 4396.87206420044, 4390.86964753769, 4343.08568737051, 
    4334.16244098773, 4318.34484114637, 4311.85174633048, 4300.56018650199, 
    4269.50039500803, 4200.25924596289, 4101.76420738588, 3972.33381563759, 
    3821.90370602495, 3687.60407449871, 3541.19410410763, 3415.98897500926, 
    3318.47402379603, 3268.1892219329, 3288.49092561094, 3387.2978515625, 
    3519.66603907519, 3688.72181216485, 3823.67404528817, 3929.50673185287, 
    3969.4684402952, 4013.38759121336, 3976.76119469723, 3896.94449739692, 
    3858.2869662973, 3848.35229690683, 3861.84676521308, 3901.48298138913, 
    3958.86746696482, 4030.96250349173, 4071.84550424681, 4092.40267864, 
    4106.70522476116, 4137.6820437937, 4150.982947172, 4180.1588662445, 
    4214.29399166683, 4246.78113513979, 4239.20635926329, 4002.5809585027, 
    3660.23683379488, 2362.87820599067, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    2922.17748475915, 3976.25673994739, 4563.48668347045, 5018.70417610578, 
    5244.92973292234, 5378.53771329888, 5476.62408950614, 5500, 5500, 5500, 
    5500, 5435.07392495528, 5277.58205174957, 5041.64644336404, 
    4809.75028521335, 4565.88356271831, 4315.20193826066, 4105.40578785493, 
    3871.39224989008, 3636.27444145827, 3361.30619888776, 3174.78655072805, 
    3144.33314163618, 3259.5328742339, 3472.82509535469, 3695.85907237597, 
    3979.74176691555, 4238.21894304981, 4419.18185522252, 4523.49535592357, 
    4536.26537701475, 4541.44240329622, 4522.92466481813, 4519.35457265469, 
    4630.06737157424, 4912.33662538795, 5167.57274188757, 5324.44685859759, 
    5320.3866761466, 5222.4460163406, 5033.66435822791, 4807.70094703564, 
    4540.85771790787, 4196.77074278091, 3671.50222142571, 2948.20526273486, 
    2092.20200493095, 1375.28154311486, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    1308.38569369017, 2093.96874809166, 2782.38026010576, 3419.21458822898, 
    3835.09358186416, 4026.26901878342, 4047.89373791036, 4047.89373791036, 
    4065.89147763595, 4174.89623571068, 4009.53422596153, 4050.25172149904, 
    4050.25172149904, 4050, 4050, 3569.65028295785, 3279.99236093096, 
    2928.1197902296, 2727.26988268419, 2514.8601470307, 2574.54700838716, 
    2875.34907384666, 3181.73602856043, 3469.78530899617, 3750.83795137173, 
    3842.87940934137, 3794.98982714292, 3662.56589503187, 3484.19605718687, 
    3323.82175924327, 3193.86342155644, 2763.34007724181, 2481.92798967904, 
    2903.56106748629, 3897.13991973993, 4645.921666684, 5090.34743792703, 
    5233.7577653576, 5259.65914915583, 5267.48858424402, 5243.6959617149,
  5124.5691318719, 5049.95965987562, 4992.04250692125, 4976.2197211455, 
    4910.78822386084, 5034.97330367623, 5022.91104306591, 4817.10156399823, 
    4483.0299200904, 3825, 4700.22423479209, 4936.72649134478, 
    5056.35300650664, 5061.61899702618, 5110.64507902312, 5076.66549167462, 
    5113.14694515635, 5113.14694515635, 5129.40062048827, 5129.40062048827, 
    5072.16075983097, 4835.63676611141, 4367.25171316883, 3501.15410150605, 
    2919.98043991929, 2058.19945217643, -0, -0, -0, -0, -0, -0, -0, -0, 260, 
    260, 543.62711826946, 750, 900.06081491837, 1608.01121097956, 
    1590.94665536754, 1828.19809706765, 2149.23494818716, 2791.67549924018, 
    3094.62727108435, 3253.26947204999, 3292.53031755643, 3364.17372019116, 
    2886.83714863844, 3007.69150315107, 2747.53049926204, 1556.63130353799, 
    1177.59008000978, 552.580141300005, 270.610395222517, 170, 70, 60, 0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 1684.35603970423, 2607.23486806238, 
    2942.40047209745, 3262.06815118504, 3988.65635192897, 3950.26284465197, 
    4039.18560125729, 3477.18717538482, 2269.62677068838, 1802.76237610016, 
    1851.63756652446, 1882.6209572581, 2027.91875165631, 2093.27317290686, 
    2222.23700167382, 2735.0062367966, 3186.92944694772, 3387.2978515625, 
    3479.5132896655, 3552.78771907862, 3638.02685221214, 3839.35064142512, 
    4160.41507504685, 4476.670277331, 4823.80501185523, 5123.50101863763, 
    5251.62964745478, 5272.13800578712, 5210.47234219571, 4948.16278816212, 
    4972.48299615449, 4864.28633422883, 5036.28057030488, 5169.96911296537, 
    5365.60990774523, 5500, 5500, 5500, 5352.61047330935, 5080.85216812409, 
    5075.99061364193, 5038.31537178516, 5041.38663054495, 5120.67395477649, 
    5028.80160770733, 4715.17465884778, 4340.52472734496, 3982.21243854093, 
    3962.57668864101, 4067.31690956173, 4115.44995165855, 4358.07320606843, 
    4842.33998136053, 5072.28359168563, 5229.93307788899, 5278.72328738851, 
    5197.11407310694, 5133.21796986305, 5043.73005220975, 4982.31755719717, 
    4849.2925811355, 4944.07500317229, 5002.50752189602, 5057.65125839474, 
    5079.72331139598, 5019.88479047043, 4878.21863704119, 4795.14066463334, 
    4649.31546763306, 4479.01490518077, 4300.42952702361, 4120.72550778431, 
    3998.52633776505, 3999.51742420088, 4126.26584032513, 4302.36653827068, 
    4433.99837933023, 4469.84727434451, 4574.20438648258, 4612.52886338224, 
    4677.9492499403, 4672.77235580333, 4623.30016393142, 4590.11110595356, 
    4545.03873192027, 4531.07942905268, 4462.13241466156, 4428.36791770306, 
    4460.14380756593, 4470.24459557349, 4385.26538093946, 4347.72657653897, 
    4330.60753472645, 4328.34015214243, 4308.55289114279, 4270.87659771475, 
    4222.76640315532, 4143.71124153518, 4050.77563134836, 3964.8653471322, 
    3834.34780984009, 3624.73774490751, 3500.82185861459, 3360.25384691009, 
    3270.27989323983, 3242.4048639956, 3323.39498290564, 3457.77640595565, 
    3623.29344234172, 3742.93796313634, 3844.98587146981, 3886.73155645744, 
    3911.35033392598, 3901.04566915657, 3822.55394895129, 3822.51451334374, 
    3841.47833663072, 3873.96376399641, 3897.59985904138, 3957.93813585577, 
    4029.70549963759, 4071.02306060454, 4073.30242023922, 4067.45263899904, 
    4095.28273243942, 4078.37257596332, 4095.12500640108, 4118.29386672429, 
    4168.89554946118, 4114.74811486708, 3960.17214247812, 3676.41837382535, 
    1754.99818839888, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 2655.38519301236, 
    3981.52477940262, 4572.87126060169, 5012.33643408941, 5226.94745726757, 
    5366.41235094262, 5452.47360014314, 5500, 5500, 5500, 5500, 
    5400.40838311701, 5248.5625673943, 5003.63017893021, 4807.61517416761, 
    4573.82907267503, 4334.26606547759, 4132.26672408099, 3936.25668620907, 
    3729.24727198519, 3512.48351788269, 3292.76736563435, 3220.50056448551, 
    3298.82312718813, 3451.83818073967, 3662.68581624326, 3992.96417052664, 
    4291.52830309192, 4466.98510211791, 4581.27247716055, 4563.39218766437, 
    4521.11435442442, 4494.82661523932, 4427.83251294601, 4397.44341811441, 
    4793.59970679538, 5103.44656144878, 5271.21803795979, 5236.21067757645, 
    5155.39038719042, 4968.64703876952, 4727.97743365156, 4437.72054486897, 
    4081.47295916373, 3545.81025216658, 2721.90652550995, 1709.77474292748, 
    917.30254714002, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 1047.17319828074, 
    1953.62558308204, 2767.74550276965, 3461.85370205082, 3904.65176452572, 
    4142.94010553067, 4235.62300857452, 4276.18832675756, 4309.34218298456, 
    4268.6170164993, 4009.53422596153, 4284.83558748531, 4212.73308622914, 
    4050, 4050, 3387.2978515625, 3055.3280307114, 2615.86299070263, 
    2560.80892738568, 2438.35449762114, 2977.46354201617, 3334.7689940575, 
    3564.71297833174, 3744.19543832454, 3895.25238238425, 3899.20413813478, 
    3820.29846277596, 3689.61093202461, 3429.58378576142, 3239.06236970504, 
    3258.50975677778, 2802.11141921495, 2084.01835198886, 2545.05146701708, 
    3793.17113535253, 4639.00712704722, 5097.13166517055, 5221.83801817871, 
    5227.19162472692, 5197.26204295803, 5195.83637306111,
  5124.93402059828, 5066.55596011761, 5002.36296934505, 5010.30183156852, 
    4967.13604925104, 5005.64752903228, 5008.9629186745, 4824.76413834144, 
    4431.46026018415, 3475, 4524.07187749797, 4887.49215388521, 
    5030.2517195219, 5023.35578045879, 5074.5060867145, 5054.12073500931, 
    5097.51111023446, 5053.03194662689, 5132.38182285946, 4976.09709086856, 
    4820.37243092442, 4633.43753687085, 3505.85736226004, 2709.62765189763, 
    2125.56651839383, 1339.9325745353, -0, -0, 0, 70, 70, 60, 60, 80, 260, 
    260, 385.417310565286, 850, 850, 1200.18100006399, 1361.37911562825, 
    1889.62897538753, 2013.53664872448, 2769.51557135009, 3114.06936348872, 
    3300.66416836323, 3483.79599229812, 3671.35250172799, 3699.17124213791, 
    3102.56356865951, 3102.56356865951, 2505.36699751192, 1436.21803989193, 
    930.374599086324, 270.610395222517, 170, 110, 70, 0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 2607.23486806238, 2698.88414167677, 3262.06815118504, 
    3950.26284465197, 3950.26284465197, 3950.26284465197, 3477.18717538482, 
    -0, 1891.86136632687, 1946.02133987619, 2159.319694633, 2077.9401405222, 
    2027.91875165631, 2369.00574661326, 2822.31722939401, 3143.24079355776, 
    3331.31999818064, 3402.12783195775, 3426.37311939089, 3425.31665805874, 
    3571.84856968712, 3839.9009502386, 4187.75360202037, 4650.47680871012, 
    5024.22711757813, 5209.39441432259, 5265.94097354922, 5212.70185951825, 
    4853.72605437092, 4899.42519008068, 5093.16172934983, 5190.41347010879, 
    5275.25868639848, 5450.37433728118, 5500, 5500, 5500, 5451.82687604573, 
    5143.41858983545, 5212.00409022812, 5224.65951442712, 5202.81969235142, 
    5246.75287616771, 5198.35801833274, 4883.57677302262, 4404.97611228157, 
    3970.94013175631, 4036.62120877573, 4330.7753245372, 4383.60436184728, 
    4615.0532601601, 4875.33067169395, 5063.05037628189, 5189.12621083908, 
    5228.25593853336, 5193.89168552044, 5096.0049297167, 5020.35187249095, 
    4982.02004699744, 4817.31259254103, 4902.82828116686, 4979.16890114279, 
    5022.76718016445, 5038.45572486902, 4962.34572622674, 4861.82504876204, 
    4747.24134492762, 4622.04672106408, 4500.60924313186, 4361.30319736834, 
    4244.12879002091, 4158.89300685536, 4117.7962860095, 4233.53287619887, 
    4361.87515737491, 4446.78650345524, 4511.57788082185, 4567.71669029237, 
    4618.79032584939, 4653.391654846, 4648.07274847391, 4642.2339827337, 
    4606.28033695174, 4592.80356727303, 4533.61695106428, 4470.69283378883, 
    4426.01378742727, 4477.14264964252, 4475.7710386291, 4419.18185522252, 
    4365.24505523702, 4341.2159551435, 4303.48439764576, 4279.67715543571, 
    4237.24758237656, 4227.76063079849, 4183.48732170684, 4102.887530277, 
    4021.51712355673, 3878.43901491377, 3684.72788546704, 3548.49814359579, 
    3400.95356065821, 3271.11455405295, 3227.29215747117, 3271.94553508785, 
    3430.79641115416, 3548.67279587657, 3675.82176015996, 3798.49015227672, 
    3814.14869468623, 3839.16577019259, 3854.66114295179, 3799.30563678774, 
    3788.57746684364, 3807.8020222168, 3849.25848728733, 3884.67022650585, 
    3944.72499252389, 3994.33790269722, 4037.76166361758, 4035.69300617354, 
    4013.80455771878, 4017.96055372947, 3998.4571271706, 4014.98006647704, 
    4035.61129647322, 4052.41880118316, 3970.41866473368, 3878.22396395879, 
    3250.25692540389, 1629.97774463681, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    2875.09364336006, 4015.6565551305, 4490.40165082037, 4929.34468292795, 
    5160.32906995383, 5322.87455138985, 5452.81679685468, 5500, 5500, 5500, 
    5497.44909797799, 5372.94548792631, 5220.00079767564, 5022.86937640191, 
    4833.08916071568, 4582.15324454809, 4419.18185522252, 4234.2217531643, 
    4017.88288151634, 3790.86854458441, 3604.74714227119, 3354.22274267024, 
    3194.65822204302, 3155.3518863711, 3409.71886585204, 3662.68581624326, 
    4026.53431972903, 4297.66309889573, 4476.57442653707, 4581.17512467755, 
    4661.23050284493, 4604.79607495571, 4517.72773412888, 4390.43875319533, 
    4298.81758211701, 4525.40503604915, 4834.65687214114, 5143.41858983545, 
    5167.36181000897, 5087.05721809004, 4893.39184195201, 4657.93810278314, 
    4364.46153147338, 3956.50067096354, 3341.10668362904, 2524.72933860262, 
    1416.94066443285, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 1013.99497014753, 
    1953.70536122821, 2735.64642180411, 3458.69920057837, 3938.52084773706, 
    4216.35501072365, 4340.40659743483, 4398.63281753065, 4442.75094421495, 
    4479.17093449159, 4195.65044760087, 4328.52096126849, 4328.52096126849, 
    3841.40753484206, 3476.02779431661, 3135.31050801247, 2765.90490531281, 
    2371.97278278599, 2244.45482914875, 2595.9629523323, 3303.85739120224, 
    3573.84598961759, 3770.94609626902, 3894.69923670917, 3968.963197457, 
    3982.06642213865, 3862.56508447148, 3689.63663161962, 3526.29698586583, 
    3292.18141076009, 3273.6313566953, 2915.4454480789, 2011.66424046617, 
    2377.28583930697, 3616.87133811645, 4577.38842722713, 5052.4359322303, 
    5192.67358688472, 5187.11271415729, 5154.12725907783, 5170.39755039666,
  5106.32727240386, 5042.82388485642, 4974.72637440828, 4966.90549451785, 
    4958.66966414618, 4997.09780559244, 4956.0504186042, 4779.07571895829, 
    4449.84116702445, 3825, 4500.63712867281, 4769.03065983916, 
    4930.43253619028, 4983.17009012326, 5016.02127803915, 5006.54907382109, 
    5028.69397214655, 5008.48721189831, 5051.28577101423, 4824.02846122149, 
    4525.44698071303, 3909.2646766453, 2926.65659298302, 2452.31045727266, 
    1697.12502302956, 0, 120, 120, 60, 70, 70, 60, 60, 80, 260, 260, 
    341.829650639455, 850, 850, 1116.42980928445, 1336.41666690083, 
    1760.82668653402, 1960.769933227, 2504.8026335501, 2817.03371978804, 
    3319.36887278651, 3568.25640945371, 3514.12973724375, 3709.92400935645, 
    3509.82241484469, 3323.13283660189, 2885.94695082506, 1534.68646627293, 
    1316.34951720624, -0, 140, 140, 70, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    1527.69956616663, 1527.69956616663, -0, -0, 3396.94879756603, 
    3918.96392909649, 3750.51423122849, 2732.73426599381, 2278.18630178498, 
    2061.90560742827, 1946.09714771335, 1946.02133987619, 1936.02767835464, 
    2070.13211372626, 2405.71031132097, 2766.26205513767, 3008.02904407981, 
    3149.53879406556, 3180.09172169356, 3220.56847707888, 3273.21191801089, 
    3387.2978515625, 3623.60382267599, 3974.7889342237, 4371.5653422445, 
    4790.71974827747, 5081.42678965777, 5183.9887000821, 5143.41858983545, 
    4996.64545098656, 4975.65294983374, 5160.01955574288, 5212.84243872138, 
    5398.0310156497, 5500, 5500, 5500, 5500, 5449.63677477636, 
    5314.98549649437, 5285.36906095313, 5281.29369759423, 5226.47152963654, 
    5290.74055241338, 5256.1014859453, 4951.82356616169, 4520.04622555118, 
    4083.63766140025, 4104.76337809715, 4290.25512515235, 4436.15520643649, 
    4701.74481181567, 4888.51639195695, 5054.47101860262, 5149.70058205427, 
    5150.50205840713, 5097.94482937772, 4991.84139367956, 4965.10354831041, 
    4920.79487847456, 4869.77019635407, 4951.34748182547, 4965.93132335534, 
    4967.83576252974, 4952.73018384372, 4860.8962037271, 4788.67889528023, 
    4693.91349577895, 4596.0896487857, 4522.68265801992, 4424.74550711832, 
    4320.21969521158, 4250.32167266241, 4241.52915431003, 4324.64155364777, 
    4419.18185522252, 4479.18846885118, 4527.61925188569, 4582.41656690836, 
    4622.1652675154, 4640.80710714069, 4644.18884329193, 4635.41208966401, 
    4599.02840483863, 4575.25583326688, 4541.13982994505, 4475.49715394829, 
    4465.958681135, 4458.22209028003, 4447.63457742715, 4419.18185522252, 
    4353.99249055481, 4317.27906632916, 4282.24953120565, 4269.7251480948, 
    4250.13244432271, 4222.08165461657, 4192.62096713765, 4142.6782993183, 
    4065.89147763595, 3939.99573811366, 3749.00549789772, 3597.44937528024, 
    3458.27439109565, 3336.29160709814, 3278.96006843125, 3269.28640074202, 
    3375.20016443263, 3477.96408476611, 3579.39540435203, 3675.56318794557, 
    3721.27612304688, 3756.3671087669, 3784.48752780292, 3768.14006552709, 
    3774.09995313735, 3792.56074398093, 3816.12375475355, 3855.22999037554, 
    3907.70008051239, 3944.34745002012, 3972.15822092044, 3966.91889454881, 
    3934.61375678041, 3925.70237610219, 3904.57550692401, 3907.63128023244, 
    3917.16357680063, 3942.93905033348, 3828.60246196863, 3672.22561394974, 
    3002.33083325109, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 3106.39034801209, 
    3939.46622839485, 4399.33039761469, 4822.25255808926, 5061.66900255407, 
    5255.94761998734, 5401.37520893438, 5488.18693099438, 5500, 
    5491.38856838496, 5438.64278578645, 5355.62153636112, 5207.38822763565, 
    5021.37420863374, 4830.73529519187, 4624.9098309824, 4431.57661430993, 
    4240.42271577029, 4045.47892365375, 3830.65915936094, 3628.79878843382, 
    3400.0365285066, 3252.09544278137, 3184.77353690137, 3388.17607353951, 
    3658.53296908088, 3973.33728933646, 4260.95203690317, 4462.30770467674, 
    4605.88809752898, 4688.40818989718, 4653.43379604364, 4549.10845646029, 
    4425.44025637791, 4360.3252977661, 4506.34651385376, 4656.99683915175, 
    4965.04349900502, 5035.21115603715, 4985.44430653035, 4827.43605336256, 
    4593.85227420182, 4281.48422019286, 3772.21481167435, 3107.90841149844, 
    2358.03389775721, 1458.27446253753, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    1150.83765438463, 1957.70788752208, 2677.5857040903, 3416.42792981397, 
    3942.5544334321, 4244.80497523563, 4424.54947205737, 4495.34204860654, 
    4537.42183424029, 4580.91928134987, 4526.39397807202, 4570.49457814698, 
    4379.48926474209, 3852.81308768995, 3133.27960515565, 2831.72123451895, 
    2392.08263821703, 2176.93482677102, 2379.01398443333, 2919.17901154923, 
    3439.63555586639, 3699.62479820827, 3872.45585855824, 3979.55522272965, 
    4009.28619511559, 4003.55027453904, 3884.00095833832, 3679.02715524761, 
    3480.21924999825, 3325.76047855969, 3247.78679771336, 2999.19211328045, 
    2487.79417609749, 2553.15327883494, 3550.91397499107, 4439.31702306223, 
    4960.60017759054, 5155.11015307058, 5154.82784357704, 5149.99006146071, 
    5143.41858983545,
  5062.03525022069, 4988.90252620041, 4878.17318945372, 4895.32647589896, 
    4909.65051939285, 4970.97896595081, 4932.97046094646, 4742.87334654256, 
    4442.71988377791, 3825, 4482.8833798664, 4717.38760333421, 
    4879.17246281929, 4939.80191664828, 4968.34691954152, 4950.44812999859, 
    4976.39365298196, 4954.39921441741, 4900.03924601299, 4622.18393288465, 
    4205.8571375405, 3241.139701056, 2470.75351147253, 2022.93259242339, -0, 
    -0, 120, 120, 60, 50, 50, 50, 50, 60, 180, 260, 330, 750, 750, -0, 
    1208.7085282568, 1553.68528288406, 1870.51785128316, 2513.22557951004, 
    3113.90056402908, 3422.8235473923, 3488.35720303488, 3368.15796448367, 
    3636.6063763028, 3511.98376184233, 3248.62961082308, 2773.24919695586, 
    1589.98416755916, 1342.42581722013, 657.807241188975, 140, 140, 70, -0, 
    -0, -0, -0, -0, -0, -0, -0, 1390.80583315737, 1558.04951571539, 
    1682.83619646607, 1782.95207135619, 1782.95207135619, -0, 
    3133.03665957874, 3131.3256583127, 2540.64680322803, 2305.37305866849, 
    1935.05359591651, 1824.24051211386, 1892.61091077732, 1882.5807990298, 
    2113.87590797692, 2368.97123300332, 2709.32519302684, 2934.31699867297, 
    3015.86712147386, 3065.78548661781, 3172.57410570258, 3239.86489802655, 
    3334.26987069889, 3526.83614073488, 3817.22448440796, 4162.99955197234, 
    4577.74968296538, 4936.70377400274, 5108.04039700166, 5097.51739499921, 
    5035.44908822513, 5120.88329095887, 5219.08625469167, 5310.7069015412, 
    5492.49924307498, 5500, 5500, 5500, 5500, 5374.89633054927, 
    5312.60370432232, 5274.84501250206, 5267.47435901498, 5236.15791963781, 
    5280.62204824533, 5297.31100552275, 5049.19699441884, 4640.29162152879, 
    4192.97027802844, 4072.88097120099, 4266.50385439167, 4539.56036856108, 
    4802.6395403807, 4935.59786863754, 5041.67254327275, 5112.36147717173, 
    5093.03141614484, 5043.81545235427, 4970.34462692604, 4940.82940631412, 
    4903.74374579262, 4939.64932194015, 4953.7678238944, 4918.33812833041, 
    4903.09778916185, 4897.34085878155, 4806.86846717799, 4732.95953506742, 
    4651.32330109995, 4582.31642897593, 4538.48294277769, 4474.22349968892, 
    4389.13494443156, 4320.68616987451, 4324.75339209082, 4379.23931642676, 
    4449.26210365097, 4495.68521063081, 4535.27148751687, 4578.94073083046, 
    4616.85557031147, 4636.28935494164, 4639.00412006492, 4625.82370664064, 
    4596.11164574604, 4568.06524834959, 4549.34294033806, 4495.94190763966, 
    4466.38646486245, 4456.57717819134, 4431.53872233817, 4381.30172268941, 
    4332.6797429472, 4294.47465045069, 4275.50129214859, 4263.18279197886, 
    4244.33152103649, 4227.004371819, 4213.30067245346, 4172.75523802854, 
    4097.91041936388, 3976.28298754407, 3814.67331352455, 3645.5751551968, 
    3506.09548126767, 3400.60474213357, 3332.56994331093, 3287.12264894429, 
    3351.92849536669, 3432.67812506059, 3503.73071602909, 3575.90165166423, 
    3644.94196549244, 3701.90019937841, 3733.91764622424, 3722.04108988203, 
    3740.79954553639, 3760.66973162685, 3785.09493162137, 3814.60883036623, 
    3858.04491751644, 3890.67867268264, 3905.43872986193, 3882.16723184379, 
    3844.26824229413, 3827.60589052005, 3801.22599352758, 3789.30998326306, 
    3790.84850348529, 3819.99745426889, 3691.15223590566, 3517.95709432001, 
    2843.67399417537, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 3183.64418214184, 
    3911.89894554823, 4338.36236357949, 4728.82048962522, 4969.04423255441, 
    5177.88436747071, 5338.20466599106, 5429.99036299777, 5453.80996873503, 
    5422.93452922553, 5380.91657721686, 5313.90953944486, 5184.65434058123, 
    5057.75743224819, 4878.24645168591, 4683.72249874214, 4491.21354142996, 
    4284.36912135024, 4077.36960158966, 3863.95694140919, 3649.28427778608, 
    3412.63107217929, 3252.52283729977, 3235.44560036547, 3418.69403026986, 
    3670.33871398812, 3953.22525591024, 4198.91670367803, 4429.11704988329, 
    4588.0816180521, 4683.54513669759, 4681.74108846227, 4603.04295262703, 
    4474.3442651309, 4371.02529356057, 4471.94150664546, 4574.56187764263, 
    4841.02567818556, 4900.37223693725, 4890.81366492575, 4758.0575137011, 
    4531.07051131776, 4182.78337648793, 3623.59818669333, 2942.29979200053, 
    2227.7092590716, 1349.42860243807, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    1147.52250999902, 1894.13449231533, 2616.02412508634, 3367.3422974446, 
    3927.74098673514, 4269.42815552544, 4475.24502554685, 4586.64771531773, 
    4640.08870406078, 4696.91864607222, 4705.17830638972, 4677.13087268338, 
    4450.5169294951, 3921.376781592, 3068.80409405792, 2619.20549226097, 
    2159.4058604481, 2088.12302146738, 2579.32542960705, 3205.24008158781, 
    3590.52205306215, 3814.14510109816, 3923.63416710136, 4038.90412822991, 
    4038.90412822991, 4019.50965194506, 3880.70098336676, 3659.22320999318, 
    3446.90378166058, 3327.72124468542, 3286.48177376014, 3147.32210416354, 
    2787.70725318521, 2745.7676376516, 3516.21952413703, 4396.82698637736, 
    4923.10180247729, 5124.12410983326, 5120.47981534954, 5116.84257605191, 
    5108.11917144466,
  4993.66163048483, 4919.55778658161, 4761.65832969925, 4797.650690221, 
    4863.39464732325, 4923.08694480026, 4891.53931575778, 4702.18248170805, 
    4395.35878581159, 3825, 4431.1981418207, 4667.61025632355, 
    4843.83372627103, 4871.81187402638, 4909.70709442532, 4908.0335509243, 
    4936.15160861974, 4879.95763664376, 4650.36391095887, 4266.25177106436, 
    3757.24426277422, 2674.2859302826, 2082.25417213134, -0, -0, -0, 40, 40, 
    40, 50, 50, 50, 50, 50, 180, 260, 330, 670, 670, -0, 1040.28651310076, 
    1040.28651310076, -0, 2781.15689994204, 3200, 3478.84204392952, 
    3423.55884688262, 3342.92841287814, 3357.11046469656, 3221.41895270135, 
    3037.5836143567, 2395.63459396248, 1593.05650296908, 1284.92450515216, 
    657.807241188975, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    1280.12060546875, 1440.88038459097, 1554.8060315441, 1656.28091056425, 
    1782.95207135619, 1870.98215458536, 2058.9427816652, 2505.62328383743, 
    2505.62328383743, 2400.3038717744, 2145.33284219989, 1820.1097607631, 
    1812.96486969767, 1897.39349779963, 1939.54486794542, 2156.88844405407, 
    2372.8767889426, 2745.65142162718, 2903.29681684049, 3000.86414129062, 
    3131.761788347, 3224.90416357374, 3271.59268718356, 3349.58615100436, 
    3478.9419892832, 3725.58598253556, 4015.76203813724, 4419.18185522252, 
    4779.07571895829, 5001.8854970266, 5008.63799229418, 4993.85702402063, 
    5127.00435321168, 5273.2109295342, 5438.29756323892, 5500, 5500, 5500, 
    5500, 5482.00825397976, 5284.95365973482, 5283.7504490526, 
    5166.37910452776, 5169.66806021184, 5251.43732455082, 5266.54779162148, 
    5319.60654642677, 5148.85504290248, 4784.15586934464, 4344.46197924365, 
    4189.81103197956, 4375.90552049447, 4663.486041781, 4897.18891172304, 
    5022.85406777496, 5097.78067621176, 5098.3505578828, 5081.86709893834, 
    5015.56145116326, 4957.33957865965, 4909.55289237953, 4890.36704906876, 
    4939.3393236299, 4910.75877507128, 4853.83972662984, 4830.67507780469, 
    4824.31077169437, 4758.53202493314, 4676.33849196111, 4626.7905699739, 
    4576.70373703826, 4542.75584876258, 4483.14596610633, 4437.50973885776, 
    4390.19147188854, 4394.93377673262, 4423.52798451952, 4483.57728127858, 
    4505.8490928635, 4541.7223941725, 4569.48398146052, 4603.20317438816, 
    4620.65272490828, 4633.68381921894, 4613.07649576746, 4598.00820840608, 
    4568.08577202072, 4544.02790648582, 4501.00480277287, 4472.68289292333, 
    4461.92420356974, 4429.26702511744, 4373.17385767465, 4321.12483168221, 
    4286.75338015639, 4273.9398189551, 4259.92999150746, 4241.26990985877, 
    4234.04073464017, 4227.5029222983, 4200.37863342671, 4127.35596779718, 
    4014.90702694158, 3875.70225877535, 3721.27612304688, 3571.87756056234, 
    3473.04237775185, 3395.58837752948, 3336.60887452732, 3358.32314853422, 
    3387.2978515625, 3439.41169983369, 3495.33133906842, 3562.07206776221, 
    3635.77139980393, 3670.42545669015, 3681.20984371493, 3695.98958768964, 
    3708.34071555613, 3728.28292320116, 3749.78130730745, 3782.7339325885, 
    3806.57266152279, 3810.44487655511, 3772.13180055759, 3728.66158333312, 
    3703.36271148403, 3667.11910684903, 3642.57880978455, 3621.18282498094, 
    3641.80868174841, 3536.89264869111, 3339.96691201413, 2707.46473650797, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 1521.67303209301, 1968.58963064644, 
    2466.81058546672, 3281.39745881421, 3850.45716064723, 4284.25597360202, 
    4626.0219964006, 4865.38155438239, 5086.71292610699, 5257.94184904955, 
    5353.74309863381, 5381.54860316977, 5361.18595849738, 5326.80186588186, 
    5279.078645203, 5167.97746758417, 5071.6089920005, 4918.65822610584, 
    4734.68087755673, 4543.41941450971, 4340.15070358661, 4112.72452563246, 
    3902.44472041344, 3675.63782302978, 3439.34712967462, 3254.53553256471, 
    3294.28158999866, 3470.82945178762, 3721.27612304688, 3982.5613996017, 
    4200.30229778748, 4419.18185522252, 4558.15168222857, 4645.09196363649, 
    4668.11964988722, 4593.63650712152, 4524.1627904442, 4438.30981538565, 
    4498.78712923443, 4596.15240115171, 4759.22234601059, 4764.28279384996, 
    4762.11704131392, 4660.40200257267, 4425.14791642072, 4024.60128199136, 
    3458.52362875294, 2817.08613874278, 2044.1318190444, 1203.40483484015, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 1103.5504492601, 1807.63017016553, 
    2553.16493236533, 3283.69742076269, 3894.25048492616, 4269.19783029536, 
    4504.88387341855, 4654.97401485086, 4732.42680196872, 4791.34115280317, 
    4827.07908413628, 4807.68871615223, 4536.39132078973, 4004.49153529396, 
    3166.91115567229, 2429.01947301561, 550, 2248.15106733755, 
    2881.30168883405, 3429.73098665546, 3759.99822320886, 3920.39564997252, 
    3983.84658323562, 4080.50538895338, 4102.95105279546, 4033.55911855607, 
    3864.15237852702, 3622.60531347122, 3399.8075592657, 3308.08139868554, 
    3366.41616407249, 3307.05538925465, 3109.81665987471, 2950.59643408772, 
    3513.04003660406, 4366.68680818266, 4866.77830460034, 5071.54757968134, 
    5070.61816960384, 5064.50130317512, 5056.9297721961,
  4947.00140112878, 4888.06508853952, 4688.28628283186, 4718.8559459201, 
    4817.51104570858, 4877.91950134883, 4848.09653287162, 4660.34784907465, 
    4332.97779351224, 3625, 4360.93774192464, 4635.60342671453, 
    4806.1837199218, 4830.8765172887, 4864.38800565485, 4861.9691443806, 
    4907.51576002365, 4768.44672489376, 4457.38288768384, 4030.43436582506, 
    3209.88030349434, 2285.41929863365, -0, -0, -0, -0, 40, 40, 40, 40, 40, 
    50, 50, 50, 50, 130, 330, 670, 670, -0, -0, -0, -0, 2820.79242438977, 
    3200, 3292.63056748436, 3292.63056748436, 3115.51086454195, 
    2933.81258394286, 2855.29103789244, 2554.50610567935, 1949.96817363022, 
    1536.75085934067, 1050.14213907029, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 1265.68394172196, 1416.07173524409, 1498.16050634527, 
    1532.65502305947, 1562.76012718202, 1679.0609863565, 1870.98215458536, 
    2058.9427816652, 2157.27970169924, 2442.04363677206, 2389.72580226072, 
    2086.98843033634, 1840.52468256066, 1836.27672348947, 1902.75109151286, 
    1993.9123264314, 2228.46542929123, 2475.0013150241, 2852.25195931826, 
    3002.30750447265, 3134.95701454803, 3280.3202603871, 3323.06829066577, 
    3350.87820114794, 3415.92727148962, 3504.08984873698, 3721.31426972542, 
    3978.15235818727, 4343.55656924247, 4661.27482700444, 4862.192374825, 
    4873.55035195622, 4966.92793397708, 5088.06247294891, 5268.66277705977, 
    5445.5885761107, 5500, 5500, 5500, 5500, 5480.70894642355, 
    5273.08345454959, 5223.73718509652, 5150.19932064213, 5107.10748918436, 
    5200.80118202288, 5260.19668323534, 5317.85634910741, 5209.89924094616, 
    4896.55771808596, 4504.0760800001, 4364.32743582896, 4573.09593944311, 
    4802.31275233026, 4961.10956836731, 5084.62103899903, 5102.95053246685, 
    5122.2578652315, 5080.74054483385, 4999.20207367216, 4908.53844669223, 
    4880.3494536835, 4905.27203324423, 4904.98960290333, 4871.73635730808, 
    4804.98393488837, 4781.32004645698, 4767.14438043069, 4724.90068552665, 
    4658.70661925141, 4617.92172152228, 4563.7684512499, 4532.34871830725, 
    4489.12492557125, 4444.25838720794, 4419.18185522252, 4419.18185522252, 
    4453.60267522763, 4497.41955207182, 4512.52851487247, 4537.22619910382, 
    4551.06725800129, 4581.48083277744, 4603.19970712093, 4621.31922447651, 
    4602.1421112027, 4589.85149475405, 4564.44698175375, 4544.46457961318, 
    4515.17523388407, 4492.84842231734, 4472.75861693691, 4434.64211662247, 
    4373.40008472078, 4328.63162307747, 4295.97015556045, 4278.04252621843, 
    4260.48313195351, 4244.76589931519, 4242.32409553101, 4234.81235649148, 
    4211.15536659203, 4142.26392730556, 4034.10336658875, 3914.24855897133, 
    3783.06982987885, 3642.5075775506, 3551.17306586798, 3474.22391088755, 
    3416.95381265102, 3389.71780375423, 3358.57140949007, 3388.01798419447, 
    3435.19854725405, 3511.40867584522, 3572.22198689742, 3614.52004290256, 
    3640.35993982091, 3650.65055782417, 3658.84349311726, 3667.7043442052, 
    3685.7068670964, 3708.16870112966, 3721.27612304688, 3721.27612304688, 
    3645.76526606968, 3582.37436937793, 3563.77916244698, 3537.7881625079, 
    3501.15230203407, 3471.14780196592, 3454.7747196652, 3359.75428544349, 
    3161.28979122253, 2582.86523506008, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    1704.93566717851, 2317.08277982653, 2758.41088867188, 3375.0151242893, 
    3759.77081088063, 4157.88507113981, 4546.0964408579, 4802.51641642613, 
    5017.37089012778, 5187.25503100212, 5287.9847172861, 5328.27544718177, 
    5317.01759772041, 5278.74632793024, 5225.79745364229, 5152.99956638484, 
    5063.8195055862, 4940.25754152749, 4779.07571895829, 4568.49207034034, 
    4379.80143999347, 4157.23888992976, 3948.55425163061, 3698.22087371987, 
    3466.76151535175, 3288.78303388005, 3332.80962335629, 3529.569628617, 
    3768.9895711114, 4015.26269115983, 4215.81921617105, 4419.18185522252, 
    4567.74855172809, 4658.50051141333, 4685.62980806771, 4594.70232343239, 
    4552.31981910804, 4460.90608045921, 4475.71933502755, 4561.10971181982, 
    4650.53528566698, 4683.33250058601, 4639.83282632802, 4545.93608241779, 
    4306.68601170722, 3857.09272759221, 3314.22175822244, 2612.73009189718, 
    1755.52698806524, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    1705.76782113248, 2500.77675879317, 3209.11722551655, 3825.26879793784, 
    4242.18003375476, 4504.28382113123, 4672.23205545649, 4780.13182041275, 
    4847.70005032461, 4901.74868261314, 4890.61637970831, 4623.06566077334, 
    4095.07981428421, 3309.76317720367, 2525.71884699404, 2231.81701066573, 
    2601.02585085934, 3198.46224440363, 3610.70805521686, 3864.35043263508, 
    3953.97839808577, 4053.46049752978, 4118.72607835438, 4128.52664222786, 
    4032.18010826648, 3844.30870751663, 3585.23142250003, 3359.85542995341, 
    3280.46915879539, 3435.68041514772, 3451.04694372371, 3366.09245597468, 
    3242.66025689234, 3583.14257694939, 4338.70836696133, 4803.11209630408, 
    5022.18542876101, 5038.26883343898, 5028.60604094739, 5015.41076607929,
  4916.06564605993, 4857.54793267947, 4650.53273673452, 4683.23949194132, 
    4779.07571895829, 4831.153446223, 4806.21332401605, 4619.5487222398, 
    4319.76945465807, 3625, 4298.88889711223, 4602.62520354981, 
    4762.57230907717, 4795.66122078171, 4818.26844875559, 4820.44457694906, 
    4846.10773503298, 4624.44742839579, 4246.42967562468, 3751.10516040804, 
    2671.41470174499, 1944.1875494432, -0, -0, -0, -0, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, -0, 330.022443918357, 620, 620, -0, -0, -0, 
    1800.82100684941, 2746.51283205854, 3352.53508895071, 3366.61213779719, 
    -0, 2347.80256219948, 2347.80256219948, 2323.32874762293, -0, 
    1341.56884446857, 1341.56884446857, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 1415.57618300235, 1415.57618300235, 1523.20169383191, 
    1533.80652121011, 1484.53527674914, 1536.52353696163, 1677.39186888901, 
    1847.32263196367, 2006.00520795844, 2076.12787160523, 2374.287939872, 
    2289.07349145846, 2070.33310971294, 1875.29560491889, 1842.86391331329, 
    1901.44151213451, 2044.1629347095, 2317.05414215977, 2611.61528153284, 
    2991.01264109571, 3194.05971724278, 3347.41810537133, 3444.75423318718, 
    3472.57964379429, 3467.40737263304, 3505.7385850753, 3570.00081844638, 
    3769.13186757787, 3993.74889813386, 4295.48757649619, 4534.62498766993, 
    4737.1375440169, 4819.33425781752, 4938.41223652747, 5047.39504672579, 
    5248.88440143807, 5416.99877737944, 5500, 5500, 5500, 5500, 
    5476.31124208315, 5250.08304305668, 5203.73794619558, 5167.62085482242, 
    5025.07308065097, 5143.41858983545, 5260.30056312614, 5312.21673513661, 
    5253.24495071545, 4975.72481624501, 4670.09800073001, 4611.70867288434, 
    4766.04112915969, 4934.60581090723, 5037.14736439613, 5129.71836065132, 
    5129.71836065132, 5128.12825174663, 5059.32320059512, 4958.7904311705, 
    4853.85297999177, 4857.20946649639, 4898.30099868081, 4872.96082650134, 
    4843.18666959867, 4790.17943847847, 4749.90458876723, 4728.68352518935, 
    4706.90951523878, 4651.06221541662, 4597.28697075516, 4544.36546266014, 
    4524.57508455402, 4487.91512724152, 4435.86995123262, 4419.18185522252, 
    4419.18185522252, 4445.69420197405, 4486.61932448783, 4499.23976264818, 
    4521.00989141526, 4529.93809153894, 4559.72050780805, 4578.29168369531, 
    4601.55396833303, 4590.22730577025, 4571.83190341052, 4549.9484462066, 
    4544.93752972538, 4530.61656141213, 4522.33326690919, 4494.93651674881, 
    4447.02870271109, 4384.50281853104, 4335.73244933652, 4300.40059996863, 
    4278.60134105819, 4260.12898959482, 4249.70511841944, 4246.13762843846, 
    4235.83332514741, 4219.62044055571, 4155.78907692635, 4050.55815241802, 
    3944.82593095239, 3840.78111980707, 3732.03903746957, 3640.88418314281, 
    3568.73301457609, 3499.76167489216, 3442.75859434237, 3387.2978515625, 
    3387.2978515625, 3388.1324371304, 3454.49614456888, 3509.10720339406, 
    3559.32537343945, 3590.65631095078, 3598.62210977812, 3608.55699422749, 
    3609.78707765383, 3619.43560315019, 3633.38551742604, 3633.79578087791, 
    3575.39368064511, 3465.12624431119, 3405.23346969953, 3395.20535790965, 
    3387.2978515625, 3346.19279419222, 3310.65529819367, 3272.01077159153, 
    3135.27148643454, 2952.43465215294, 2468.01522134192, 230, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 1697.12502302956, 2065.17916448128, 2643.1261766284, 
    3065.78548661781, 3512.78671827774, 3843.42798382039, 4178.91912772059, 
    4495.36221648255, 4746.06066082042, 4949.74941407975, 5102.08270913917, 
    5197.80259985708, 5252.86001240995, 5241.87366979274, 5197.09981787791, 
    5149.94453368945, 5125.00308172207, 5050.24156564761, 4928.05245363938, 
    4779.07571895829, 4578.39783902876, 4391.18127572491, 4186.03969655444, 
    3978.31330538147, 3725.38033356872, 3500.98518382071, 3321.3232664705, 
    3387.2978515625, 3598.36053641957, 3834.38641265388, 4051.14985849122, 
    4248.83522409485, 4448.31321228436, 4600.79572421334, 4696.998328222, 
    4735.50704117915, 4661.08229454579, 4581.85105858686, 4466.02170987524, 
    4432.75501647491, 4481.65388635622, 4553.83927888484, 4545.26769755156, 
    4516.84356448207, 4408.34223533659, 4140.58393452371, 3696.72831745299, 
    3092.7823512614, 2291.23626524634, 1503.99728863726, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 1597.38097966531, 2437.51962075667, 
    3117.40598876986, 3705.41176157014, 4177.71820636248, 4475.04700732103, 
    4672.67254940881, 4799.7307913782, 4880.29935694982, 4940.76926669186, 
    4938.58846180915, 4706.21875476103, 4221.72261407297, 3531.57960300106, 
    2933.66681531184, 2690.43337824479, 3041.1411746906, 3480.9664973067, 
    3806.17060738757, 3969.44567411953, 4032.00950024784, 4143.44169004707, 
    4166.66866400854, 4159.61338097924, 4036.57326584705, 3821.94633897536, 
    3549.10609329575, 3333.90756648808, 3252.60955077267, 3491.92572064955, 
    3584.68645643142, 3542.19468583443, 3471.78134439951, 3664.16985306492, 
    4311.16472939041, 4740.80976806014, 4967.72856562793, 5005.40348089866, 
    4995.69064325307, 4993.30234720702,
  4889.26420288856, 4817.0463201364, 4618.93166848822, 4644.23033390462, 
    4731.3129960573, 4763.85673035034, 4763.85673035034, 4581.4368682588, 
    4307.06166739764, 3625, 4256.23390071616, 4558.33198755672, 
    4722.17765300654, 4765.28086609869, 4779.07571895829, 4781.8798475681, 
    4740.75541549945, 4453.43405033939, 4018.33347911251, 3345.09753581579, 
    2269.17880281278, 1641.84320407244, -0, -0, -0, -0, -0, 40, 40, 40, 40, 
    40, -0, -0, -0, -0, 370.154968261719, 550, 550, -0, -0, -0, 
    1717.76242473643, 2727.11091376977, 3200.3661237562, 3235.92035697326, 
    2676.03421139656, 850, -0, -0, 1044.78738711101, 1044.78738711101, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 1815.87238679557, 1815.87238679557, 
    1656.20056807915, 1576.5176349341, 1500.00413948834, 1508.36507136229, 
    1665.75933220759, 1820.3121269146, 1910.44413469881, 1990.26323416523, 
    2173.84404209685, 2441.17646957166, 2287.51174502973, 2097.10422791177, 
    1905.07548894355, 1836.78054626628, 1935.05359591651, 2118.94836689101, 
    2438.29983931444, 2758.41088867188, 3161.42357319319, 3394.85154736976, 
    3579.89936585396, 3634.18101743251, 3637.95984082378, 3618.53696960508, 
    3613.88678998521, 3664.73637820108, 3838.71687555794, 4021.57023645501, 
    4260.10995829635, 4444.5522441601, 4639.81049525209, 4779.07571895829, 
    4884.7890273905, 5044.88726765572, 5238.73832165219, 5391.84768159519, 
    5490.59071244554, 5500, 5500, 5500, 5437.19555978395, 5279.85760735382, 
    5213.42603638524, 5166.22314453637, 4969.43508046709, 5143.41858983545, 
    5274.69192712983, 5320.25791178552, 5279.1260289044, 5070.31625317266, 
    4842.35380730899, 4829.6879124229, 4921.48423007799, 5045.44663564866, 
    5106.83741797193, 5161.37937607366, 5151.92599795408, 5116.53938813569, 
    5029.31878864086, 4927.75928812731, 4820.78791271194, 4839.13880827302, 
    4872.39930518123, 4841.35935348269, 4813.89302046708, 4767.90644594144, 
    4730.46391444583, 4700.5555153572, 4675.10351717003, 4624.35715918169, 
    4573.13515719694, 4531.68730034221, 4509.55329144353, 4478.14108658737, 
    4434.30533595579, 4409.16991235783, 4399.90735668768, 4423.02792368045, 
    4457.81948165381, 4475.78561577237, 4497.98060944656, 4509.55422834723, 
    4534.74122286319, 4541.77868924111, 4573.04634418613, 4575.17850459951, 
    4556.33424623948, 4533.12105568411, 4543.11155559041, 4544.23698623764, 
    4547.07653616627, 4520.94750879879, 4463.75493269124, 4400.62428209927, 
    4339.24313676789, 4298.98759448811, 4273.79408521532, 4258.25845975424, 
    4249.78917324482, 4244.4261701137, 4235.33140112133, 4224.74264820034, 
    4165.58808899849, 4068.61271604436, 3971.36725941413, 3877.56068978074, 
    3793.72353207274, 3721.27612304688, 3647.22719236298, 3568.09301717835, 
    3495.6326205727, 3426.656165121, 3391.52484482185, 3359.01662060654, 
    3405.45561755699, 3458.59124294368, 3509.5962543933, 3537.32486810292, 
    3545.59490322127, 3554.47180595575, 3552.27045746992, 3554.54384959498, 
    3559.47132634212, 3523.43816874922, 3395.48762564442, 3251.79066076327, 
    3190.28151517521, 3194.20516812796, 3195.96012837159, 3179.3360923988, 
    3147.27833820404, 3093.95590081846, 2938.47819242442, 2740.07923563202, 
    2367.22827460219, 230, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 1760.93870041925, 
    2022.62921130954, 2466.66776221529, 2945.32057855141, 3306.00313955129, 
    3669.99021852421, 3960.9336299952, 4244.95727713257, 4467.56973624438, 
    4689.15227490468, 4871.59256196043, 4998.19318187208, 5087.21725627025, 
    5131.68388122042, 5122.40585954291, 5076.21079778062, 5046.56320346766, 
    5065.69241380102, 5014.62823268397, 4911.19568956749, 4779.07571895829, 
    4585.72752090394, 4381.05567637462, 4181.58513956013, 3982.42235220299, 
    3743.25481779995, 3531.725193756, 3387.2978515625, 3448.04207501048, 
    3677.12297545958, 3913.55686966446, 4106.55631253271, 4306.36761458443, 
    4492.05357305678, 4654.99281109757, 4748.61526057677, 4748.61526057677, 
    4733.48905749933, 4638.85534485255, 4507.8103288903, 4419.52481283243, 
    4427.44182061166, 4444.62063306743, 4434.94204621657, 4383.37678301496, 
    4240.86350942333, 3943.06171637988, 3492.86907956938, 2817.78873060332, 
    1956.79605494691, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    1499.48238589581, 2362.16572511306, 3027.87940237769, 3573.30072449102, 
    4086.10957417187, 4419.18185522252, 4653.23394173825, 4800.04510077447, 
    4897.77116230154, 4965.21761841694, 4970.43043613092, 4798.83163338095, 
    4382.70797050461, 3794.96617516495, 3359.64966075422, 3162.98821904907, 
    3432.3949654237, 3738.93985173426, 3995.09390567723, 4086.34520858216, 
    4144.32084551644, 4239.85655697625, 4235.34250022944, 4184.04777268771, 
    4035.44152924804, 3789.00280369041, 3523.8637503017, 3309.76983006846, 
    3253.72716016327, 3522.77983878495, 3669.70561515102, 3654.2574544338, 
    3584.71332779515, 3689.53837420734, 4246.85513832929, 4674.61243729438, 
    4909.49781716254, 4969.87214142747, 4959.47490142524, 4963.73513778312,
  4860.83175673281, 4779.32003499337, 4611.41293582602, 4632.19583199269, 
    4706.61574961338, 4755.77176934146, 4729.29157785071, 4540.50208047838, 
    4285.13914886571, 3625, 4239.05327649845, 4515.85155559564, 
    4687.58741497443, 4739.81148967958, 4731.02204384531, 4742.97047558393, 
    4651.53224586341, 4325.44145923465, 3809.06850897817, 2913.60193880017, 
    2033.68151658251, 1538.53108067165, -0, -0, -0, -0, -0, 40, 40, 40, 0, 0, 
    -0, -0, -0, -0, 405.889248404243, 1525, 1525, -0, -0, -0, 
    1743.07338488654, 2617.36454292325, 3017.62213576729, 3032.84207394675, 
    2676.03421139656, 2356.13889038631, -0, -0, 1044.78738711101, 
    1044.78738711101, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    2049.20051658534, 2049.20051658534, 1784.22437651528, 1603.32605539082, 
    1484.00331440451, 1574.18337977744, 1802.25010200423, 1910.84580190342, 
    1975.65294105126, 2126.67494623239, 2401.62947105329, 2401.62947105329, 
    2389.68812353883, 2144.21275112439, 1922.75427224132, 1852.01181951735, 
    1974.88600480617, 2200.35164434631, 2552.29233586565, 2875.3074386521, 
    3312.63852293163, 3582.86894848281, 3757.5845512409, 3791.02617059697, 
    3785.53736301248, 3732.37373184769, 3702.42926410957, 3763.7797200265, 
    3914.26430389488, 4065.89147763595, 4236.10539420052, 4401.11402492975, 
    4581.86055992574, 4661.26930460831, 4780.37658215922, 5038.29874074687, 
    5238.45656679924, 5379.52824326193, 5463.04690286548, 5500, 5500, 
    5492.48048731205, 5383.72848241374, 5283.48706976107, 5218.58351169914, 
    5182.78398300401, 5031.74737897957, 5160.98753893228, 5268.52248140026, 
    5332.33661863774, 5303.90921765153, 5163.9551122162, 4985.72585034129, 
    4965.25281460548, 5024.36931788783, 5109.80610557133, 5156.20342863862, 
    5180.39354783935, 5155.08334656732, 5099.10793709106, 5007.08649634825, 
    4901.6229039107, 4810.83010129434, 4815.54964864406, 4835.07366068643, 
    4806.97258177085, 4788.65628562071, 4745.97432646592, 4714.34777897668, 
    4678.05118237265, 4645.90354571641, 4598.09365794181, 4551.41385945408, 
    4512.94916580832, 4491.43815279276, 4467.59692910188, 4431.2423995165, 
    4403.58172823507, 4385.68792855562, 4403.37885256657, 4428.96980682514, 
    4453.97888115922, 4471.79702480049, 4486.80279487443, 4506.49370219169, 
    4510.8033393009, 4545.025168037, 4557.73327071599, 4539.96065760023, 
    4522.34741370624, 4535.96891441904, 4551.76183317607, 4560.01064252199, 
    4540.99218253621, 4478.19471895355, 4419.18185522252, 4346.90761862552, 
    4297.1316327739, 4269.23566046013, 4253.30192530734, 4245.36943925461, 
    4235.98046901504, 4230.05938502757, 4225.80203641345, 4171.98868530167, 
    4081.97029398452, 3989.19966216198, 3897.69153105027, 3824.86572567133, 
    3755.56881037207, 3692.38183532531, 3612.18470053863, 3536.27268724208, 
    3462.69103628593, 3396.96973275101, 3341.87764169758, 3375.78631207792, 
    3423.15729101994, 3471.70886049689, 3493.3967007436, 3501.30510250751, 
    3504.52304942477, 3502.55137109305, 3502.98394829963, 3494.78483441442, 
    3408.43598803512, 3236.27389823937, 3074.99206445468, 2995.12195692016, 
    3011.17933124086, 3049.90596883012, 3050.65640621809, 3019.96783315914, 
    2943.10276560037, 2788.92235995439, 2597.22168680332, 2260.92851362099, 
    230, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 1923.01065577414, 2373.92968654752, 2796.28485232837, 
    3178.79854165604, 3465.58006532342, 3794.25776153109, 4071.89323646863, 
    4290.61573370208, 4454.78395625412, 4643.37019658836, 4801.90534987497, 
    4902.42949748358, 4980.47663072119, 5009.74588035331, 4996.30574029975, 
    4962.20678459009, 4946.97365025329, 4983.3294662939, 4969.64989986326, 
    4880.18819186686, 4726.6368638155, 4551.7572848737, 4365.7990491059, 
    4158.49120391624, 3963.22595993371, 3754.02464291806, 3548.78794948776, 
    3433.80112547313, 3515.62055995909, 3743.0211432822, 3974.8010192818, 
    4176.08621391638, 4373.81290991437, 4547.73610095671, 4710.08287042092, 
    4792.02662364736, 4824.13113602507, 4790.7247573797, 4698.36057566346, 
    4567.50207242202, 4458.56719104606, 4408.94729011916, 4363.55092307675, 
    4348.32181328712, 4255.94954384883, 4094.09279768155, 3764.18709272835, 
    3294.86525292472, 2575.39376681714, 1755.5000883053, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 1424.2878185178, 2253.04416431318, 
    2942.33148026134, 3475.26762050009, 3993.91845607336, 4364.34670342382, 
    4625.27699015553, 4788.26724364775, 4899.88902194131, 4971.4838868374, 
    4984.33752267145, 4850.65765465894, 4501.59711196152, 4004.05164716144, 
    3685.13476203639, 3519.82545917055, 3698.13522745452, 3921.87935757841, 
    4129.50069099641, 4196.49823806352, 4243.87154227552, 4313.23588045686, 
    4291.77148430532, 4208.2613727918, 4027.17749916758, 3752.29456162268, 
    3500.8498535364, 3300.14351703175, 3281.81555968497, 3546.66406946059, 
    3695.6563606193, 3695.6563606193, 3605.43598203457, 3659.22260334288, 
    4187.5321303631, 4599.52528839763, 4859.19938374804, 4933.96046996008, 
    4936.46444284118, 4937.24165710596,
  4836.69061075695, 4744.67464145838, 4615.51740931935, 4634.3907992737, 
    4684.01140242921, 4727.00388015416, 4693.34577937498, 4505.58187911926, 
    4266.42190056547, 3625, 4230.69342137927, 4488.21181386812, 
    4657.91973588695, 4704.73448195399, 4683.48741193616, 4694.75561238142, 
    4520.57634708076, 4184.90479661589, 3542.09294487648, 2477.71130359074, 
    1806.22866574856, -0, -0, -0, -0, -0, -0, 40, 40, 40, -0, -0, -0, -0, -0, 
    -0, 405.889248404243, 1675, 1675, -0, -0, -0, 1679.83710582827, 
    2339.44884540419, 2743.33277354079, 2731.60748061094, 2559.76854293381, 
    2277.96407951909, 550, 683.282409667969, 844.978224970989, 
    844.978224970989, -0, -0, -0, -0, -0, -0, -0, -0, 2436.22417775844, 
    2678.80829523527, 2604.90809910833, 2215.65191696498, 1861.60324905306, 
    1670.4240340854, 1550.44297987013, 1677.42764473313, 1961.32641827885, 
    2067.47636420707, 2111.62276085452, 2441.7417010315, 2723.61175040764, 
    2723.61175040764, 2564.79222526643, 2192.68514354182, 1943.0511526816, 
    1877.98755690185, 2032.9690974491, 2295.68690941253, 2680.84965824862, 
    3015.1661047121, 3483.2903973121, 3775.00339382627, 3920.70381830304, 
    3960.04064660614, 3934.34962166974, 3845.72564798857, 3807.50040954474, 
    3879.38687119163, 4009.92129110006, 4108.33704566865, 4218.2785668845, 
    4374.40566644351, 4512.7333216722, 4537.82362159089, 4695.12617865027, 
    5009.61504186288, 5226.92367078828, 5376.38231916787, 5439.94791750142, 
    5500, 5500, 5447.57033481051, 5310.40240872951, 5257.62249408015, 
    5230.9883874909, 5203.66638040503, 5151.58136001077, 5203.5152767624, 
    5276.65121486721, 5339.20574177692, 5341.94126867427, 5254.40687398641, 
    5105.87938659928, 5080.88873027691, 5103.7338394324, 5179.70406617473, 
    5202.53100737671, 5184.4023606421, 5143.41858983545, 5068.34852309324, 
    4973.78310052548, 4853.40258718535, 4789.07514413498, 4779.07571895829, 
    4784.73241936018, 4779.07571895829, 4753.63050140858, 4717.72478817635, 
    4687.49966943258, 4654.20844534993, 4616.40112376786, 4566.36719957925, 
    4517.25473903687, 4490.70210924306, 4466.90178897321, 4448.93790745146, 
    4419.18185522252, 4392.65233798394, 4365.97128343537, 4383.43499613415, 
    4398.59455294315, 4427.05294882329, 4433.91075570778, 4455.66731040104, 
    4465.04464892016, 4483.4099738166, 4516.00589906264, 4533.97986689636, 
    4518.67574286219, 4513.36196908498, 4529.18197708674, 4553.61671645264, 
    4572.11413640666, 4557.06593676871, 4492.78804503797, 4426.97150255388, 
    4353.95652009705, 4295.25545689192, 4264.95064266963, 4241.88238453149, 
    4238.05621165792, 4221.73167764427, 4219.24735104942, 4223.83928703492, 
    4171.14301158905, 4090.77632060877, 4005.08914616779, 3917.35190889549, 
    3850.47008991175, 3784.81183040405, 3727.80596543668, 3653.52972084628, 
    3575.78422169938, 3485.57034689121, 3397.1525600772, 3327.53541622011, 
    3350.3422276539, 3389.59095950051, 3432.35128059052, 3446.76025408762, 
    3452.04402335411, 3450.80993443621, 3448.40572158328, 3448.97462607877, 
    3418.80657852862, 3287.37934854641, 3077.35396457073, 2885.96724362981, 
    2786.40049501772, 2821.59726882768, 2892.0242388402, 2922.54994793205, 
    2879.2086532369, 2779.88735971922, 2627.01888124141, 2430.57346253498, 
    2169.94576218929, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 1312.12389170436, 1725.56190095196, 
    1974.04001948795, 2263.62873339504, 2715.72999644099, 3101.46442879662, 
    3409.04895765303, 3657.61005376247, 3951.34357010608, 4178.6207359668, 
    4327.8124683909, 4453.35797286401, 4599.44282046924, 4726.77040484657, 
    4791.18827340132, 4847.54324156549, 4850.84342569185, 4834.6266569701, 
    4800.19828045835, 4808.67037593659, 4861.70843464308, 4868.78899913043, 
    4809.31764804645, 4650.60591930772, 4479.68709098923, 4331.2322368523, 
    4127.2894897248, 3933.0884738908, 3762.5212328676, 3571.33253223163, 
    3492.52164154939, 3606.70505565176, 3820.46425021694, 4053.74971226621, 
    4263.7720491925, 4459.84542644615, 4625.00014330782, 4779.27482194878, 
    4849.42039014939, 4864.22055633635, 4833.55073644407, 4744.38641470878, 
    4618.27007636741, 4512.60623804472, 4405.06777279459, 4315.23902209634, 
    4240.6840761949, 4127.13741687097, 3917.71986794557, 3558.95099947741, 
    3088.8037044564, 2339.12447644165, 1597.65565434226, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 1309.13904996341, 2098.50962011158, 
    2835.55398309637, 3387.2978515625, 3867.44269601395, 4293.79208848563, 
    4582.25901248047, 4763.83542212402, 4884.94992711522, 4973.0133834084, 
    4998.4290079395, 4900.11277008008, 4640.21557606358, 4245.0996094361, 
    3955.8070919045, 3810.72436020261, 3961.34284877521, 4137.62443977769, 
    4271.87398634701, 4303.14785907224, 4335.98249293, 4376.40734838024, 
    4344.98026900543, 4234.62962395179, 4029.4145515682, 3726.40418994299, 
    3483.68747677087, 3290.30393478131, 3310.3344412651, 3582.83236861736, 
    3798.19261359347, 3726.83688225287, 3606.47397479246, 3595.07040664511, 
    4113.43611080294, 4509.55314525094, 4797.33989828286, 4894.34963505849, 
    4912.41974366457, 4909.78685263187,
  4815.72193956269, 4732.4877764652, 4618.54807290123, 4648.38703814551, 
    4670.71624764866, 4700.44593679683, 4664.43454307983, 4487.01358457205, 
    4290.99801875003, 3625, 4317.78716937001, 4503.72597497363, 
    4629.03793972681, 4674.68083780318, 4645.40388958995, 4613.81972235165, 
    4430.93331660149, 4120.69414246182, 3222.47120404996, 1855.2425573029, 
    1443.69849303831, -0, -0, -0, -0, -0, 40, 40, 40, 40, -0, -0, -0, -0, -0, 
    -0, 376.184461505711, 1875, 1875, -0, -0, -0, 1315.78797400763, 
    1559.24280407439, 1977.93417332144, 2060.11381577896, 2119.53861839732, 
    1967.8170014119, 550, 683.282409667969, 683.282409667969, 
    664.235845920315, -0, -0, 892.753383279219, 892.753383279219, -0, -0, -0, 
    2346.66404046463, 2868.1452132177, 2868.1452132177, 2768.13939054295, 
    2304.30552694, 1815.02528472016, 1706.90759175403, 1538.72280125643, 
    1659.93613597978, 1936.9619604055, 2141.88797015525, 2295.05356095948, 
    2711.35059732483, 2728.57603304067, 2728.57603304067, 2686.31523294629, 
    2205.76225372227, 1935.05359591651, 1885.38529340538, 2077.26805113516, 
    2366.92270644395, 2835.53135740642, 3102.81778860575, 3660.39544446101, 
    3930.06650274095, 4100.66611694744, 4137.18442953292, 4036.22543583118, 
    3940.51044836923, 3879.69695522245, 3998.49094349275, 4118.34477400734, 
    4125.27622610855, 4242.23870338991, 4377.15518214207, 4374.40566644351, 
    4242.1594229728, 4756.04471906385, 5007.01528845477, 5246.04274134923, 
    5374.39469748172, 5409.30982198879, 5462.97805881767, 5445.5472700677, 
    5433.63804442417, 5223.18966112854, 5115.40903031512, 5267.48748887493, 
    5236.81983204715, 5287.56451389306, 5258.48134812842, 5269.97698392817, 
    5327.03876230401, 5401.72643489933, 5292.92165545496, 5205.669523982, 
    5165.9827220174, 5185.86671759594, 5226.96758515395, 5234.60364770671, 
    5174.61913869916, 5106.98241769903, 5038.39940313714, 4937.83175631361, 
    4746.56583951835, 4741.51255836311, 4722.58579343065, 4760.2199229661, 
    4744.03670392015, 4729.60646952939, 4703.75889878034, 4678.60637012881, 
    4642.78824880801, 4580.31651695464, 4521.53713433229, 4482.69074434152, 
    4455.79494114558, 4437.01864069736, 4425.24915170715, 4382.91638918628, 
    4380.4659597342, 4340.02249716903, 4359.32603858139, 4387.31459808471, 
    4399.86580705686, 4419.18185522252, 4439.64004417288, 4430.01686989184, 
    4456.49232560226, 4484.29739018186, 4504.93059263896, 4499.45200975234, 
    4490.40780879219, 4520.59676364085, 4559.65627632647, 4588.07385222532, 
    4580.77138979406, 4512.91160594137, 4444.21175359692, 4359.93986113336, 
    4286.69401991833, 4256.39908600929, 4235.65294675013, 4238.15408638195, 
    4199.05546420313, 4193.91845200409, 4227.94352057658, 4176.8390121132, 
    4095.31623509756, 4028.32697564577, 3936.05711574249, 3870.46988968638, 
    3809.91590885199, 3759.79093673808, 3688.1397551329, 3606.86312259996, 
    3504.84384962875, 3389.862006339, 3295.11554422499, 3330.54927481829, 
    3366.23763683526, 3397.23329574831, 3408.81861251097, 3405.29272440325, 
    3403.05308542135, 3396.87624093911, 3401.12411482542, 3331.65673622809, 
    3196.39684768435, 2961.80215697572, 2758.41088867188, 2614.34221212947, 
    2663.37420250981, 2763.680348037, 2794.60831831274, 2703.52703186401, 
    2586.08990919284, 2401.69604566808, 2265.72683500488, 2152.21274431087, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, -0, -0, -0, -0, 
    495.553629324057, 880.898309915524, 1518.09675270997, 2081.66625245757, 
    2361.6373615267, 2761.3452990267, 2964.72426890236, 3335.28167508886, 
    3627.86839083239, 3899.80010521169, 4117.70944226277, 4273.23621888103, 
    4375.98997004855, 4464.04464621472, 4563.80196458022, 4666.21567044031, 
    4708.82177282505, 4725.55034841535, 4714.29690842642, 4668.1956454847, 
    4575.58078059113, 4597.97149999138, 4690.28081276694, 4738.61590210354, 
    4675.12713683385, 4570.00648483904, 4364.81435090758, 4247.25198287839, 
    4099.56172433861, 3933.66832060753, 3748.23918341874, 3585.40467200259, 
    3555.98090715257, 3698.65961880288, 3900.04656833852, 4158.30856826067, 
    4337.51696627623, 4540.9460314527, 4707.91711671645, 4861.25072853061, 
    4937.22757482151, 4924.72967355532, 4895.28773867949, 4779.07571895829, 
    4657.45254223999, 4549.40277323586, 4361.25673422925, 4256.01666904329, 
    4173.68820587389, 4003.90750907539, 3734.95570833335, 3319.92791374239, 
    2941.1191673571, 2027.94697249728, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 1679.47715043407, 2728.26635183864, 3293.40365138752, 
    3758.03617193986, 4228.30112126213, 4546.85102623334, 4740.61020595747, 
    4869.58314957633, 4966.44205376598, 5015.81755186656, 4953.3249157716, 
    4791.43871123542, 4419.18185522252, 4215.36513284437, 4120.093416686, 
    4204.43216572402, 4306.3009284202, 4377.39199200627, 4368.08840350501, 
    4422.30095224566, 4448.46214372164, 4421.95126022169, 4253.95784613598, 
    4008.57634651079, 3761.80247572479, 3482.12217403858, 3218.45303220371, 
    3296.77567338721, 3619.23491864801, 3849.26063739397, 3770.81602760998, 
    3593.78137076092, 3410.18761140455, 4065.89147763595, 4420.81072004438, 
    4743.29481232435, 4868.97584346368, 4891.19314267991, 4892.51639324417,
  4795.29509895905, 4721.72194771532, 4641.80774720683, 4635.42502800344, 
    4640.19395319281, 4666.5136660734, 4629.33425337513, 4501.24472258633, 
    4239.32274645323, 3828.56570930226, 4266.70375389599, 4456.78300050944, 
    4594.32275274774, 4636.81784483265, 4629.94190666417, 4586.45176234573, 
    4233.80894122256, 4003.06261239173, 2573.80838383234, 1850.5848196105, 
    1058.40966742668, -0, -0, -0, 0, 40, 40, 40, 40, 40, -0, -0, -0, -0, -0, 
    -0, -0, 2075, 2075, -0, -0, -0, 550, 550, 0, 1350, 1350, -0, 550, 
    661.526418862301, 661.526418862301, 661.526418862301, -0, -0, 
    1228.73264249509, 1310.30091507123, 1416.37009771951, 1723.2482264083, 
    2137.39733164616, 3146.67760393543, 3065.78548661781, 3119.60562841953, 
    2987.4708654721, 2423.58839083251, 1920.32646721917, 2078.82192465023, 
    1990.90474292726, 2103.09221850126, 2266.0172869958, 2339.97434845484, 
    2800.5701523625, 3365.6029227297, 3365.6029227297, 3096.76360166797, 
    2808.42200508649, 2278.70600200967, 1990.8759066269, 1944.42126957376, 
    2123.00198998638, 2437.72126289661, 2927.82837693857, 3298.25476867872, 
    3801.48769189991, 4071.05528986661, 4217.8258988056, 4210.29245731329, 
    4143.20950201397, 4005.18469422313, 4002.09172027912, 4088.86093467206, 
    4188.12446713097, 4195.27849200386, 4260.74763527819, 4376.55810240604, 
    4207.71612039642, 4471.64792609743, 4465.80094786992, 5130.21712275631, 
    5261.34910817823, 5369.09823877868, 5344.61248088066, 5401.45771515803, 
    5375.91682018484, 5363.08521992117, 5171.66986125905, 5170.36363698645, 
    5294.31864909627, 5301.52438930354, 5322.25725494246, 5331.52904909389, 
    5323.94041957056, 5334.29805174819, 5339.54860787582, 5256.7771255343, 
    5239.00195954472, 5218.89557645897, 5218.13230987805, 5230.37222846335, 
    5201.47883093758, 5164.85973270428, 5000.84118707779, 4963.47355136227, 
    4810.9975741715, 4697.62816486953, 4550.46650531267, 4696.90112406717, 
    4731.76196302689, 4709.75208276565, 4710.0316834496, 4667.61587552193, 
    4646.65013726124, 4620.25652753683, 4540.73646153282, 4456.36513110911, 
    4419.18185522252, 4419.18185522252, 4403.73359500317, 4404.83141146798, 
    4383.25150473393, 4369.48484852888, 4344.15811955713, 4337.80431937772, 
    4336.57658218167, 4364.56418218347, 4383.94495714227, 4403.67161123652, 
    4400.89710034319, 4442.38024195805, 4455.56341320709, 4496.61744445455, 
    4489.86093302932, 4473.24598583792, 4516.18023528396, 4564.00805860021, 
    4583.77770603462, 4582.73851600792, 4513.91524865686, 4446.70114435439, 
    4360.24616780477, 4290.22313702265, 4230.79646118611, 4218.14464124783, 
    4212.01206599467, 4190.08518842975, 4179.91350950121, 4208.26623552173, 
    4161.90403791061, 4083.68868846915, 4020.14476255031, 3923.60005867064, 
    3868.21272493129, 3810.36155411672, 3757.63841129152, 3704.81399532351, 
    3624.72587454762, 3525.44706863354, 3395.96424625048, 3301.12745817507, 
    3303.23023524112, 3342.16363152921, 3365.66487115253, 3376.96859037819, 
    3365.41641064838, 3369.77372285449, 3364.03012873379, 3363.54185830651, 
    3284.86089796966, 3103.62266389669, 2862.18405958349, 2286.30936547391, 
    2113.85456139861, 2267.39830311673, 2514.4872721108, 2621.92081881528, 
    2614.25881653879, 2441.94107249612, 2262.1389531927, 2105.45741664448, 
    2064.07911294137, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 0, 658.013178042496, 1116.72772899215, 2195.07758275949, 
    2642.89099152197, 2998.40755552941, 3167.10906680034, 3174.20816640038, 
    3505.82017695958, 3887.06079898086, 4045.93739071162, 4192.68007044086, 
    4324.84437796705, 4353.3942017092, 4426.87490715916, 4487.55769432059, 
    4534.24763181948, 4480.4132390598, 4519.25443809027, 4466.6014992956, 
    4483.81358629141, 4421.74760835457, 4479.46731392532, 4590.52210557589, 
    4614.89794215313, 4599.78782706719, 4500.3763879064, 4306.8939580823, 
    4114.33308207284, 4019.59300645207, 3927.12427995501, 3789.01311747851, 
    3588.24082023025, 3640.7091691621, 3796.56788345808, 3994.51463740077, 
    4190.43824049261, 4427.96857494485, 4587.62839753961, 4780.15361069728, 
    4900.95470664607, 4963.34388513065, 4970.90852167764, 4927.45560773195, 
    4817.93109757465, 4680.1392236943, 4550.86499200533, 4419.18185522252, 
    4290.45693824512, 4137.29685518299, 3890.42480294228, 3444.2900677012, 
    3242.23384884989, 2758.41088867188, 1732.46260674385, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 1385.42172725573, 2480.47589069406, 
    3144.62441895564, 3627.10837386603, 4120.49809941976, 4485.28428871354, 
    4697.49639426882, 4847.90277054832, 4953.20340825618, 5016.13579492634, 
    4983.12059796919, 4859.67400563373, 4564.94235167895, 4404.08750975959, 
    4303.44081312716, 4320.41955333929, 4382.75259013627, 4452.7425453771, 
    4425.78718219212, 4473.16324413113, 4466.10288489181, 4433.36958993963, 
    4268.92759924942, 4039.02736435581, 3777.36156089927, 3473.82482577941, 
    3225.15887399638, 3309.62204746803, 3605.61345980866, 3810.28117892563, 
    3810.81773267156, 3536.87892912011, 3278.24191286381, 3924.33337526522, 
    4362.86067596739, 4672.79398079188, 4822.04590702735, 4854.45128923295, 
    4859.95690669978,
  4750.02511212146, 4687.18326632177, 4628.69380212755, 4612.11171134758, 
    4606.61591079491, 4641.18561888279, 4601.0428166663, 4446.81479312492, 
    4192.98608298982, 3893.9638109611, 4225, 4395.24316057961, 
    4565.62970974935, 4599.85461820868, 4602.43102503245, 4501.56866921556, 
    4121.02312588949, 3605.92348226993, 2418.89646089749, 1779.34859112181, 
    -0, -0, -0, -0, 0, 40, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, 2075, 
    2075, 2075, 0, 0, -0, 1587.77571008475, 2039.71855592823, 
    2158.21133074781, 2123.72584689912, 1560.07541661515, 360, 
    924.663409229888, 858.535857424203, -0, -0, -0, 1801.67026252769, 
    1788.20419036853, 2039.50703359144, 2478.51839579046, 2952.26890370315, 
    3203.03237673986, 3139.5558394632, 3097.0152544098, 2979.69321962768, 
    2727.28947462346, 2391.65874431132, 2356.56761970502, 2364.58581457844, 
    2476.60186268267, 2667.96748395476, 2965.05202607916, 3401.83231852729, 
    3660.05684695161, 3621.87603438816, 3308.26856251556, 2881.11215999562, 
    2361.40342388498, 2078.74299982884, 2027.86191551998, 2193.07195167356, 
    2497.8241502954, 2935.37385917587, 3419.43096544049, 3856.55482136552, 
    4127.37850659097, 4251.73666769152, 4249.09623033138, 4171.46024579038, 
    4081.97662625481, 4085.24983208039, 4114.05863904554, 4209.53644956827, 
    4226.55718140955, 4247.2709613053, 4299.54257742116, 4206.75139827964, 
    4518.56355790328, 4744.54889442246, 5105.72036095872, 5273.08601425765, 
    5362.80442571885, 5365.92358709256, 5363.60299040055, 5347.49208591733, 
    5308.65437600964, 5251.45887495843, 5271.5645552169, 5318.17179589295, 
    5341.72949864961, 5348.43258563472, 5347.97531812999, 5355.12782532053, 
    5377.91283734397, 5311.26003410393, 5259.81559743349, 5247.80559064118, 
    5221.7880670486, 5215.20971443686, 5211.38087726134, 5181.85766137999, 
    5125.33232011233, 5006.75628810018, 4874.39743808812, 4710.47638896207, 
    4599.35442128728, 4583.03953062385, 4633.47504007002, 4672.46295430405, 
    4672.85376457976, 4639.45757195988, 4597.62870745379, 4589.61263299545, 
    4555.20902264298, 4481.2402902453, 4419.18185522252, 4387.31356400356, 
    4392.6194588507, 4396.25171768427, 4402.65009493067, 4390.75668253264, 
    4364.48573185582, 4330.75968463766, 4328.15141500079, 4329.75386446021, 
    4348.33724665657, 4365.78954095509, 4372.45532268072, 4379.16190841631, 
    4406.14952548916, 4440.09470016689, 4468.73975245675, 4482.04492387345, 
    4489.87192886754, 4516.06016649294, 4556.60065617053, 4580.01696442281, 
    4572.41809127812, 4516.67981568402, 4438.58917343773, 4352.97207839579, 
    4277.52631984159, 4220.27875880894, 4193.37672474321, 4178.27773014892, 
    4167.61778966574, 4165.54657448113, 4165.73566248651, 4130.83823257646, 
    4065.89147763595, 3991.43349268945, 3917.34596877693, 3858.12539109924, 
    3798.75180749784, 3752.49359411356, 3701.34672931402, 3628.4966581906, 
    3521.28980544816, 3405.54740647316, 3314.93943648452, 3302.52920105611, 
    3323.69106185184, 3348.94610256262, 3356.63224634424, 3344.52929597962, 
    3345.87080881633, 3339.44736533266, 3325.48648688334, 3214.0083312381, 
    2968.36431916096, 2544.14721217489, 2074.19078561389, 1984.34252873361, 
    2151.89580297244, 2381.92698702114, 2550.76200301117, 2593.24701318957, 
    2150, 2150, 2124.41880962616, 1962.89792043278, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 80, 140, 978.799393179614, 
    1610.88941883635, 2398.11801019572, 2859.49342245896, 3165.77420906344, 
    3349.62681020471, 3518.6088629284, 3760.5972774837, 4017.31643871248, 
    4163.39039072121, 4255.90910028397, 4302.72796665006, 4313.88730376988, 
    4328.49987975982, 4322.76017070891, 4303.76025660833, 4284.10509702636, 
    4263.40286437953, 4218.14579190604, 4196.65577477688, 4186.42538186475, 
    4286.55154716921, 4427.98698336661, 4544.2078132666, 4536.06777613174, 
    4496.62679054746, 4316.73930913556, 4127.55876679028, 3969.89249757619, 
    3850.7079620353, 3824.35303336107, 3753.69564027686, 3771.29835092276, 
    3906.56404958623, 4078.46948934786, 4281.07728965277, 4460.56709283086, 
    4648.39543415729, 4820.95535332722, 4933.8311401256, 4994.87375955116, 
    5006.00165125196, 4956.46410365911, 4867.42806914463, 4742.45131625731, 
    4594.41329809079, 4456.3969080535, 4293.87334212202, 4116.86798185159, 
    3862.55924588893, 3537.29433217147, 3119.38878730892, 2598.85437924789, 
    1809.2114913985, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 2295.04015802337, 3018.38572532335, 3482.73229676571, 
    3942.65785248641, 4375.44763986092, 4643.02996668519, 4812.79424278399, 
    4935.83751030265, 5009.02664025428, 4993.05796168726, 4888.02822326973, 
    4663.79069806591, 4505.92018426188, 4401.02593194318, 4419.18185522252, 
    4451.72346798025, 4491.03239748587, 4482.5194812168, 4479.8357905396, 
    4460.33111679628, 4398.93599449876, 4253.09512071207, 4038.40856157102, 
    3746.36198608355, 3452.45878195794, 3256.31126909471, 3356.25136668615, 
    3619.99143072028, 3798.4786719666, 3740.63104468037, 3463.72617997329, 
    3258.33382727186, 3721.27612304688, 4221.54611303745, 4605.2356969386, 
    4779.07571895829, 4810.29092524396, 4805.81687257376,
  4717.20578565867, 4670.01287193038, 4610.21204811432, 4593.21511003383, 
    4588.83859719884, 4615.3626638642, 4573.1950027722, 4427.78001215648, 
    4178.34840555561, 3852.64904164094, 4225, 4357.7994714375, 
    4536.26714981535, 4572.24991666389, 4579.88888795815, 4426.4310604406, 
    4016.56112117272, 3430.20680736734, 2147.45079569013, 1607.89975560785, 
    -0, -0, -0, -0, 40, 40, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, 2175, 
    2175, 2175, 0, 0, -0, 1571.7764885476, 2098.14181333472, 
    2115.42316698416, 2069.64957443011, 1485.70309610736, 360, 
    924.663409229888, 858.535857424203, -0, -0, -0, 1788.20419036853, 
    1788.20419036853, 2397.62758126254, 2860.52812700922, 3242.13414917075, 
    3314.95752700516, 3202.27796448812, 3145.79336391937, 3081.44303623487, 
    2902.15435560079, 2681.03978433427, 2613.53315599251, 2645.82845991683, 
    2783.05673914933, 2998.74551186749, 3358.46914524402, 3765.07451066519, 
    3931.99077054955, 3765.58505591468, 3454.12666747514, 2933.78837407435, 
    2403.74423783514, 2131.52420079009, 2082.3736773403, 2241.48570669301, 
    2556.664187993, 2985.36483997957, 3506.0538167986, 3934.85012111949, 
    4192.71428502235, 4294.45863617311, 4286.85519766734, 4207.40598071566, 
    4129.99330192874, 4144.56625970358, 4157.45221519829, 4248.91885823439, 
    4240.12906390389, 4254.74492152341, 4275.58222377716, 4160.12823741668, 
    4578.0530220098, 4807.34038910863, 5121.62248324646, 5286.11314858407, 
    5364.95562364291, 5357.27222401537, 5339.81681935991, 5321.12254135563, 
    5275.18291977275, 5278.60345460995, 5301.10479106946, 5353.93771034653, 
    5388.73895764085, 5377.04033031262, 5371.88935529429, 5389.97710402816, 
    5384.09406156233, 5294.78398276195, 5250.16126174158, 5244.74617443147, 
    5224.14401057215, 5209.71356030065, 5197.3259086319, 5158.55442325542, 
    5079.52240396587, 4970.01321297085, 4795.79352395522, 4633.56803878966, 
    4520.93879219961, 4524.37648084134, 4591.46571519612, 4638.83335609884, 
    4637.17115354713, 4584.89395495504, 4546.35550793778, 4550.06757083625, 
    4516.01166414778, 4440.24902988896, 4372.26727266432, 4360.28228696346, 
    4375.70549006914, 4387.36579247926, 4399.01439013691, 4390.02353006023, 
    4361.6187682628, 4322.95898488791, 4320.26638343056, 4320.3020973032, 
    4335.10863480272, 4349.72338956765, 4350.32437766557, 4358.702020566, 
    4382.85624092161, 4421.83959091977, 4453.854190137, 4473.02197554875, 
    4489.57891400373, 4515.09717132112, 4553.71392729044, 4579.15570831318, 
    4572.6371327703, 4518.66500427572, 4439.41038899217, 4349.66862811539, 
    4269.50965450151, 4207.23294004273, 4175.44188251397, 4156.78543696632, 
    4146.47217387135, 4144.33982132047, 4140.59630711028, 4111.10238171397, 
    4045.7980068337, 3971.51693271679, 3902.0492740202, 3845.36807115213, 
    3785.95970284303, 3745.14164674024, 3699.82100754724, 3630.42950005738, 
    3521.84893113695, 3407.8710085725, 3312.22782224282, 3296.77653068252, 
    3312.57506257616, 3334.26159668588, 3338.32727493676, 3324.12654998905, 
    3321.35657932933, 3312.34224927194, 3292.22898635501, 3157.02631308476, 
    2894.14961886732, 2358.38043182363, 1870.6157436193, 1841.94758599898, 
    2054.81568342569, 2307.49672991601, 2507.21592001922, 2590.92313353939, 
    2517.01588986904, 1915, 2148.83675413454, 1972.91520646831, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 80, 140, 
    978.799393179614, 1888.78556876643, 2614.23165658547, 3074.07715228271, 
    3339.55444617672, 3533.83183365641, 3704.3410198977, 3948.69825733804, 
    4141.73571191396, 4238.32807391874, 4284.63022555077, 4301.76264468138, 
    4284.95878903042, 4254.7153934546, 4213.98532625967, 4160.32972370892, 
    4135.98871870116, 4085.50299698683, 4031.92037243048, 4008.48030260276, 
    4007.81986867346, 4145.16799063009, 4320.22780876239, 4472.91123043968, 
    4492.80557795051, 4486.96656901794, 4317.8847173445, 4118.1716131078, 
    3938.56855626755, 3827.89141510251, 3868.58356620469, 3848.34070273355, 
    3870.97556876132, 4006.90533408315, 4164.58620679666, 4355.78419090407, 
    4503.45380500297, 4701.5184560711, 4866.82378902305, 4966.95595235825, 
    5025.28253239017, 5037.14694034705, 4992.64941892912, 4907.682706136, 
    4787.8464046581, 4632.32318810759, 4473.07462264089, 4299.0968762062, 
    4097.63136060543, 3833.65765064988, 3500.13496332418, 3031.42956142545, 
    2529.88480845287, 1712.76593826216, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 2124.94664566325, 2871.35985283265, 
    3387.2978515625, 3850.43578105538, 4271.97411182033, 4596.82062431056, 
    4784.14914008786, 4925.80886125837, 5007.38690888327, 5010.47598212561, 
    4931.81722012504, 4734.50528210306, 4589.54789945688, 4401.02593194318, 
    4477.68015298619, 4499.29836655212, 4527.80116143832, 4519.07170788734, 
    4499.84098482141, 4467.37018979318, 4387.3339705486, 4237.03354833218, 
    4032.85323940633, 3726.66284560376, 3443.43386021, 3260.5524318876, 
    3376.58430559119, 3640.80562945173, 3802.06625727124, 3721.27612304688, 
    3401.09716046982, 3133.64920831336, 3597.73410133403, 4136.52837658356, 
    4545.69486921402, 4727.70839954359, 4779.07571895829, 4779.07571895829,
  4686.7, 4641, 4583.8, 4571.3, 4569.6, 4583.4, 4542.8, 4388.3, 4201.7, 
    4038.8, 4225, 4318.2, 4498.4, 4546.4, 4529.4, 4317.5, 3891.3, 3117.7, 
    1844.5, 1280.12060546875, -0, -0, -0, 0, 40, 40, 40, 40, 40, -0, -0, -0, 
    -0, -0, -0, -0, -0, 2275, 2275, 2275, 0, 980, 980, 1379.86463460185, 
    2098.14181333472, 2098.14181333472, 2069.64957443011, -0, 550, 
    557.411143006913, 140, 140, -0, 2021.36629750456, 2179.24860719026, 
    878.52111686723, 3309.18510022601, 3521.84615464773, 3521.84615464773, 
    3549.16756284828, 3243.4016174843, 3243.4016174843, 3359.43717808935, 
    3277.11828380242, 2964.5, 2912.4, 2996.4, 3168, 3387.2978515625, 3672.9, 
    3981.6, 3981.6, 3902.2, 3519.5, 2941.8, 2435.2, 2178, 2143.2, 2296.7, 
    2613.1, 3041.3, 3554.9, 3980.9, 4222.9, 4311.9, 4299.6, 4233.5, 4173.3, 
    4184.6, 4212.9, 4271.3, 4252.9, 4236.3, 4180.4, 4243.8, 4609.7, 4856.1, 
    5143.41845703125, 5308.8, 5365.2, 5347.6, 5325, 5305.4, 5243.8, 5276.4, 
    5319.1, 5375.7, 5500, 5412.3, 5398.9, 5500, 5371.9, 5290.4, 5244.7, 
    5216.1, 5186.5, 5178.4, 5170.4, 5127.2, 5038.1, 4893.9, 4689.6, 4509.6, 
    4440.4, 4482.4, 4575.3, 4616.1, 4583.1, 4510.7, 4491.9, 4506.6, 4484, 
    4423.2, 4371, 4359, 4365.8, 4380.9, 4390.02353006023, 4390.02353006023, 
    4357, 4324.5, 4319.7, 4318.2, 4330.7, 4334.8, 4316.7, 4347.9, 4373.7, 
    4408.7, 4443.9, 4466.3, 4486, 4510.1, 4548.6, 4574.3, 4570.9, 4515.6, 
    4436.9, 4348.3, 4262.8, 4193.2, 4161.7, 4136.3, 4121.9, 4111.4, 4103.7, 
    4079.6, 4021.6, 3951.4, 3881, 3825.9, 3771.2, 3733.2, 3690.6, 3626.1, 
    3520.3, 3407, 3310.7, 3291, 3304.3, 3319.3, 3320, 3301.1, 3292.4, 3275.2, 
    3246.9, 3090.1, 2810.2, 2256.5, 1397.8, 1383.5, 2075.4, 2341.2, 2544.1, 
    2641.5, 2611.2, 2262.8, 2244.9, 2040.5, 140, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 40, 40, 80, 120, 315, 2207.6, 2840, 3235.1, 3486, 
    3686.6, 3873.3, 4065.89135742188, 4199.3, 4271.4, 4290.9, 4279.1, 4230.7, 
    4170.2, 4100.5, 4052.1, 4024.8, 3964.8, 3871.2, 3851.4, 3884.4, 
    4065.89135742188, 4244.5, 4419.181640625, 4470, 4459.5, 4368.5, 4186.2, 
    3981.2, 3886.2, 3934.8, 3943.8, 3999, 4124.1, 4266.1, 4436.3, 4574.2, 
    4764.4, 4898.1, 4988.9, 5044.4, 5051.2, 5015, 4937.8, 4823.9, 4666.7, 
    4496.1, 4308, 4100.6, 3819.2, 3460.2, 2911.4, 2490.1, 1738.9, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 326.990295410156, 2696.5, 
    3257.8, 3731.4, 4132.8, 4512.2, 4738, 4896.6, 5000.4, 5018.3, 4958.5, 
    4794.6, 4650.1, 4446.1, 4504.1, 4526.8, 4549.5, 4542.7, 4507.6, 4447.8, 
    4343.3, 4202.2, 3976.7, 3696.1, 3420.5, 3285.8, 3433.3, 3672.1, 3691, 
    3691, 3329.4, 1630.02973949383, 3468, 4020.1, 4464.5, 4675.8, 4731.8, 
    4736.9,
  4656.21810608508, 4612.02991333705, 4557.46983263699, 4549.34915141438, 
    4550.2835465171, 4551.43847432756, 4512.37613167791, 4348.79947011804, 
    4225, 4225, 4225, 4278.68677955117, 4460.46545544002, 4520.61690448997, 
    4478.96316106897, 4208.63355874644, 3766.03872094921, 2805.2590095437, 
    1541.49676846218, 950.03786035807, -0, -0, -0, -0, 40, 40, 40, 40, 40, 
    -0, -0, -0, -0, -0, -0, -0, -0, 2275, 2345, 2345, 0, 980, 
    1460.05715569835, 1852.26994328192, 2181.66272587343, 2043.81592535395, 
    1955.48655624773, 0, 550, 550, 550, 220, 2578.76862955457, 
    2822.80253293689, 2856.19122074871, 3023.49917473008, 3309.18510022601, 
    3521.84615464773, 3571.1287964192, 3434.90074609786, 3308.27220500819, 
    3251.55883527115, 3206.02665542384, 3198.74870994342, 3248.00030192507, 
    3211.20626355831, 3347.01355753106, 3552.94934236399, 3761.45432562552, 
    3987.42967230866, 4198.04221514563, 4224.45844343196, 4038.77437901378, 
    3584.81012767599, 2949.82432977971, 2466.66776221529, 2224.38834896258, 
    2204.07581016557, 2351.82394121619, 2669.45762067577, 3097.32048904498, 
    3603.69609588789, 4026.92700297697, 4253.15228309053, 4329.39189826616, 
    4312.38531277147, 4259.58030191638, 4216.67731200962, 4224.55416879842, 
    4268.41688091017, 4293.60627476796, 4265.6864035827, 4217.81823916358, 
    4085.15016945752, 4327.43412080012, 4641.25045425476, 4904.90425857945, 
    5165.18849922349, 5331.41663196526, 5365.46010635253, 5337.97357685786, 
    5310.12082174755, 5289.6246855461, 5212.50642444087, 5274.143157853, 
    5337.11491868185, 5397.36828821037, 5461.98997727664, 5447.52745938488, 
    5425.91786686679, 5399.22652998864, 5359.71391283143, 5286.03191630244, 
    5239.22745252536, 5187.48137734775, 5148.76506483369, 5147.04544033366, 
    5143.41858983545, 5095.8643035663, 4996.68841591578, 4817.72836026478, 
    4583.47981725254, 4385.61752140457, 4359.93733573712, 4440.48026419224, 
    4559.07912533716, 4593.41200110292, 4529.11729314291, 4436.56942201421, 
    4437.38302155236, 4463.14801907893, 4451.99576078707, 4406.23315466667, 
    4369.7049310585, 4357.73187008085, 4355.80896263721, 4374.5082116583, 
    4389.99504927991, 4377.80459490054, 4352.46683356885, 4325.9701806664, 
    4319.15205114534, 4316.03210075186, 4326.37463990587, 4319.7834135815, 
    4283.00407448378, 4337.09509014109, 4364.54629955761, 4395.62253979666, 
    4433.95725262888, 4459.65644960819, 4482.48456331177, 4505.18746735886, 
    4543.49315184804, 4569.44212403229, 4569.20451762751, 4512.45064433307, 
    4434.35316228579, 4346.87362516287, 4256.04193611014, 4179.23205984738, 
    4147.9179558677, 4115.81027930074, 4097.40447054389, 4078.45673523896, 
    4066.86851802602, 4048.18264179217, 3997.47086468149, 3931.28788328457, 
    3859.89400129958, 3806.35307559426, 3756.36899425257, 3721.27612304688, 
    3681.29397869425, 3621.80911417567, 3518.73726750411, 3406.05487808995, 
    3309.23305311937, 3285.30566248274, 3296.00869525902, 3304.26674672988, 
    3301.69300454507, 3278.10026252819, 3263.46655704274, 3238.10810538564, 
    3201.65358538302, 3023.10813321609, 2726.17813502466, 2154.56349361485, 
    925, 925, 2096.0752046555, 2374.92114543932, 2581.02251095747, 
    2692.03743650688, 2705.39139498616, 2610.52583883355, 2340.86993911353, 
    2108.14961840607, 1697.12502302956, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 40, 40, 70, 90, 150, 1018.42469309895, 1637.71937638688, 
    2526.34770431844, 3065.78548661781, 3396.07222884053, 3632.44238589135, 
    3839.41225204499, 4042.19330166314, 4180.89564481771, 4256.93338488505, 
    4304.51487182002, 4297.25406320893, 4256.3593491048, 4176.40694443346, 
    4085.63389672371, 3987.10656065449, 3943.81314594605, 3913.518539923, 
    3844.15310620153, 3710.56082708059, 3694.33309071749, 3760.96911321549, 
    3982.18206804715, 4168.72702699816, 4359.2648891749, 4447.24488543494, 
    4432.00547682558, 4419.18185522252, 4254.21734350229, 4023.86047012171, 
    3944.54512311657, 4001.00850869157, 4039.34114238342, 4127.07818334049, 
    4241.30749720313, 4367.57254074239, 4516.72646095187, 4644.95652225001, 
    4827.27921781122, 4929.33554409994, 5010.82455168241, 5063.55697860376, 
    5065.31316496835, 5037.29781907942, 4967.92600211475, 4859.98031737742, 
    4701.01115172184, 4519.11761644024, 4316.80944049183, 4103.61409569789, 
    3804.80949875182, 3420.21711044476, 2791.45035853576, 2450.29222577449, 
    1764.99870487861, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 2521.67595412861, 3128.39104757317, 3612.2753434716, 
    3993.61626470275, 4427.49216408496, 4691.94777984859, 4867.3500999786, 
    4993.3646464327, 5026.08552626011, 4985.08705209187, 4854.63281979171, 
    4710.64658574435, 4491.23118635742, 4530.57438465511, 4554.34775295171, 
    4571.1770323065, 4566.41888686638, 4515.45203661713, 4428.32123921296, 
    4299.20069976576, 4167.39195560899, 3920.54704488982, 3665.49449080577, 
    3397.57065785239, 3311.1428222522, 3490.08483977421, 3703.42126423253, 
    3703.42126423253, 3660.80264411147, 3257.69962229477, 2929.40272862134, 
    3338.29824585666, 3903.5896808633, 4383.20935975095, 4623.8261312693, 
    4684.54828194615, 4694.76409216572,
  4621.97571487104, 4585.35956691425, 4529.56870412715, 4520.69874886416, 
    4528.89393048776, 4522.11549190925, 4487.32562298225, 4320.18429974264, 
    4225, 4225, 4225, 4238.70050485668, 4419.18185522252, 4486.25704035608, 
    4380.43761597288, 4082.04855603029, 3637.68630537534, 2578.58419796008, 
    1541.49676846218, 950.03786035807, -0, -0, -0, 0, 40, 40, 40, 40, 40, -0, 
    -0, -0, -0, -0, -0, -0, -0, 1017.10544838444, 2345, 2345, -0, 980, 
    1460.05715569835, 1852.26994328192, 2172.8015458317, 2031.87316486225, 
    1905.9833156242, 0, 550, 550, 550, 220, 2896.68611093377, 
    3137.98355699975, 3173.21045708954, 3360.23434720917, 3563.06308622327, 
    3687.62351752852, 3641.90079460461, 3501.15704458939, 3346.99104899029, 
    3318.81359308291, 3267.56619362597, 3281.41708618247, 3402.74717208597, 
    3436.47059258804, 3616.85787799547, 3813.90357251954, 4014.00533675946, 
    3987.42967230866, 4356.79351112357, 4352.54346833765, 4110.97962559836, 
    3626.46430903605, 2977.32033292094, 2512.42785034036, 2266.89417870146, 
    2257.35759496732, 2401.19244117407, 2718.17825280639, 3133.09308498211, 
    3631.79307180207, 4041.7336586352, 4262.05133198956, 4330.93203503805, 
    4317.8953482842, 4277.73219586152, 4241.34325152988, 4243.87233786146, 
    4289.14380976468, 4294.9404677489, 4257.45686307914, 4193.92767517134, 
    4049.17841231427, 4361.85391812887, 4648.50916537342, 4933.20401010244, 
    5211.71319043102, 5346.28854390964, 5375.35114783058, 5337.18405453915, 
    5302.19970964235, 5283.28989086729, 5205.72622566604, 5281.84222270844, 
    5346.95803576076, 5408.1181280465, 5482.82716510905, 5461.65305146993, 
    5445.13792282107, 5397.77540817084, 5356.677565012, 5290.09814633983, 
    5237.32816464599, 5174.8192350523, 5102.30881004275, 5110.68655080662, 
    5107.81442858785, 5065.93746072326, 4941.54884389859, 4732.50227471482, 
    4494.39971586244, 4291.15407358991, 4285.45083973661, 4419.18185522252, 
    4546.7545051848, 4569.96381227456, 4487.17406839483, 4398.95543976855, 
    4419.18185522252, 4448.31769343407, 4445.36853154215, 4406.92823526775, 
    4373.07996342842, 4362.34476722602, 4356.85013544019, 4371.5403529879, 
    4386.17235192568, 4375.39190251956, 4352.13617053461, 4328.40257636428, 
    4319.93230486055, 4318.97228217111, 4329.9907294584, 4313.53458227119, 
    4277.48839013042, 4332.13241595209, 4358.40285106393, 4389.45290570025, 
    4427.28395961115, 4453.58594898469, 4477.15502316646, 4499.9133574134, 
    4538.07781864005, 4562.33912162714, 4565.26988248946, 4506.71342208664, 
    4435.12938388763, 4348.68062564532, 4255.89863929078, 4175.68755568415, 
    4134.10507295422, 4100.53182106772, 4072.88425154998, 4048.0645253683, 
    4038.0677577591, 4019.1951755695, 3972.90151299347, 3914.33677183027, 
    3844.5092958164, 3789.97937991733, 3741.05199480054, 3706.91386550914, 
    3671.1804751546, 3615.43245962153, 3515.074111675, 3406.79740345728, 
    3306.59688092324, 3280.23410425679, 3288.88908825705, 3293.29896718128, 
    3286.15130295593, 3258.67812819556, 3231.58639770788, 3204.55450464482, 
    3152.3729817352, 2963.26514913148, 2674.10920679691, 2168.52280430137, 
    1050, 1924.98723006532, 2117.06455765732, 2397.84031136778, 
    2605.95683973695, 2738.97452000469, 2738.97452000469, 2703.79724816451, 
    2493.46392439911, 2244.19556874557, 1808.11386874274, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 40, 40, 70, 150, 150, 1018.42469309895, 
    1959.77203072735, 2803.49095686921, 3293.42352469521, 3620.46290369599, 
    3809.73145613214, 3981.00877621936, 4142.63117046521, 4234.11089562674, 
    4282.55904123062, 4290.24474287073, 4266.284021928, 4200.63976652775, 
    4095.45206563412, 3974.97334041478, 3869.08701492765, 3826.70271864143, 
    3803.38874839623, 3754.49586864116, 3710.56082708059, 3694.33309071749, 
    3721.27612304688, 3927.76427579, 4127.21590973158, 4350.73303984822, 
    4461.88308034403, 4459.49345468124, 4460.68683669596, 4312.76836751356, 
    4023.86047012171, 4034.90951909064, 4094.4577564559, 4126.22936073289, 
    4222.25017017035, 4329.68698268315, 4449.23207383725, 4576.33364685625, 
    4709.13728870396, 4864.25575305454, 4956.37750358789, 5021.4066302044, 
    5069.93948447285, 5073.577395048, 5046.65847881389, 4982.92484446581, 
    4880.4976458725, 4722.81749671946, 4538.62490553224, 4330.28243089235, 
    4110.94237122556, 3796.33823720444, 3399.6972938097, 2736.28595423963, 
    2435.43030157465, 1804.5058854672, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 2333.12530434629, 2958.22235702567, 
    3486.30453697816, 3908.89446147116, 4313.37331404613, 4636.99641905176, 
    4840.71872302143, 4984.55375988535, 5033.33191519258, 5006.73244710615, 
    4889.72414455217, 4747.01706401228, 4519.08254437327, 4539.71703172546, 
    4571.84352564569, 4578.54063362494, 4568.44274102337, 4507.90666779309, 
    4401.01916229676, 4260.48342933137, 4117.62115231287, 3866.03573942457, 
    3639.19585417013, 3398.24334956257, 3332.76462594204, 3506.85923075774, 
    3732.65369390538, 3832.74929566191, 3630.84136725168, 3205.88069313824, 
    2833.94457824672, 3234.44489415736, 3805.41839001912, 4287.57531436188, 
    4567.79744846136, 4644.46488533637, 4655.11286844402,
  4583.2, 4553, 4506.3, 4493, 4497.9, 4490.3, 4455.8, 4289, 4187.5, 4187.5, 
    4187.5, 4192.3, 4373.6, 4373.6, 4260.8, 3925.6, 3468.2, 1245.9305357383, 
    200, -0, -0, -0, -0, 0, 40, 40, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, 
    -0, 550, 2550, 2550, -0, -0, -0, -0, 604.567051525335, 1905.9833156242, 
    1905.9833156242, -0, 180, 894.244117986666, 1562.20971658541, 
    2242.99485598024, 3315.23597617876, 3529.91562028298, 3577.83281210703, 
    3813.83476969017, 3883.6869272165, 3883.6869272165, 3841.98086450999, 
    3338.93057922864, 3299.91541073171, 3242.31901984739, 3293.8, 3401.8, 
    3579.6, 3666, 3843.7, 3997.7, 4192, 4227.4, 4488.8, 4445.9, 4138.5, 
    3635.4, 3014.5, 2568.9, 2332.3, 2322.5, 2473, 2774, 3175.1, 3656.9, 4044, 
    4260.2, 4326.2, 4316, 4283.6, 4264.9, 4257.9, 4304.9, 4268.4, 4230.1, 
    4142.5, 4074.8, 4376.1, 4656.9, 4968.4, 5234.8, 5366.2, 5388.5, 5325.1, 
    5294.3, 5269, 5194.2, 5292.6, 5353.6, 5419.8, 5500, 5500, 5500, 5402.5, 
    5352.9, 5292.1, 5242.1, 5182.7, 5109.1, 5097.7, 5070.9, 5016.7, 4868.7, 
    4629.2, 4364, 4198.9, 4231.6, 4406.3, 4532.6, 4537.4, 4468.6, 4399, 
    4423.3, 4458.1, 4462.9, 4425.1, 4391.1, 4381.5, 4365.6, 4373.4, 4383.8, 
    4379.1, 4358.6, 4334.7, 4320.1, 4323.7, 4335.3, 4323.2, 4299.4, 4337.7, 
    4354, 4385.3, 4423.2, 4451.5, 4472.8, 4495.1, 4532.7, 4559.6, 4562.5, 
    4508, 4441.4, 4355.4, 4267, 4183, 4126.8, 4085.5, 4051.6, 4023.2, 4009.8, 
    3987.6, 3949, 3896.5, 3830.9, 3775.9, 3731.2, 3698.1, 3660.6, 3604.1, 
    3509.4, 3405.3, 3308.6, 3277.4, 3288.7, 3295.9, 3281.3, 3241.2, 3210.4, 
    3174.4, 3095.8, 2901.7, 2617.6, 2191.85375976562, 1312.5, 1952.4, 2139.4, 
    2404.8, 2615, 2768.1, 2820.3, 2802.9, 2625.9, 2401.2, 2040.1, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 0, 60, 90, 150, 150, 1478.68884277344, 
    2339.6, 3080, 3530.4, 3806.5, 3963.2, 4089.1, 4200.5, 4256.6, 4269.7, 
    4240.7, 4190.8, 4109, 3960.4, 3827.7, 3721.27612304688, 3683.8, 3699.5, 
    3697.8, 3681.4, 3680, 3732.3, 3942.2, 4143.5, 4354.7, 4489.3, 4537.6, 
    4541.7, 4420.7, 4211.4, 4161.5, 4176, 4224.9, 4329.1, 4404.5, 4497.7, 
    4615.4, 4745.9, 4880.3, 4961.6, 5017.8, 5061.7, 5063.8, 5043.3, 4991.8, 
    4889.8, 4727.3, 4548.2, 4331.6, 4108.7, 3773.5, 3372.7, 2758.41088867188, 
    2381.4, 1841.8, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 588.311954109153, 2736.8, 3323.1, 3770.5, 4189.9, 4547.9, 4792.1, 
    4963.9, 5031.6, 5020.2, 4925.3, 4785.9, 4590.2, 4523.1, 4581.9, 4579.5, 
    4558.3, 4485, 4366.3, 4208.7, 4038.3, 3803.3, 3586.6, 3387.2978515625, 
    3350.7, 3542.8, 3754.4, 3841.6, 3611.9, 3129.4, 2737.4, 3112.2, 3697.8, 
    4193.6, 4485.3, 4581.8, 4602.7,
  4544.40413647167, 4520.65045317626, 4482.9912161561, 4465.38511327129, 
    4466.90680460461, 4458.56381711997, 4424.23589191163, 4257.72513729267, 
    4150, 4150, 4150, 4145.92493353926, 4328.01451152459, 4349.86461609365, 
    4141.26154998286, 3769.23019980531, 3298.61842894775, -0, -0, -0, -0, -0, 
    0, 40, 40, 40, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, 2550, 
    2550, 2264.31309766387, -0, 2329.22323764764, 2308.180178707, -0, 1520, 
    1520, -0, -0, 1903.15576311494, 2368.03567067594, 2785.33135542628, 
    3315.23597617876, 3529.91562028298, 3577.83281210703, 3813.83476969017, 
    3883.6869272165, 3929.93672984637, 3886.99011666037, 3727.73926687976, 
    3521.25754961837, 3341.1130012539, 3319.98860550204, 3522.26408297398, 
    3756.45306780234, 3895.53081366613, 4070.44262914048, 4181.47624672693, 
    4370.07967675398, 4467.28115905241, 4620.78671968057, 4539.34235242765, 
    4166.08682348273, 3644.25932298759, 3051.74445211101, 2625.46263286592, 
    2397.72171741362, 2387.5524185162, 2544.8473590112, 2829.81794256174, 
    3217.059019403, 3682.05703110127, 4046.31708655561, 4258.3362360673, 
    4321.38452355031, 4314.18589741457, 4289.44843619805, 4288.41762854695, 
    4271.84251294387, 4320.6881540069, 4241.90627155034, 4202.79481732475, 
    4091.00986730682, 4100.48198026923, 4390.33167298487, 4665.37586653399, 
    5003.55095129469, 5257.81774780841, 5386.05933752358, 5401.71444507068, 
    5313.00879859205, 5286.48264136695, 5254.70072484264, 5182.76894318574, 
    5303.34453854377, 5360.14323471802, 5431.48145788039, 5468.2840099432, 
    5458.24677731872, 5443.71777936979, 5407.25565503018, 5349.0291767429, 
    5294.15203686587, 5246.94327486525, 5190.5342761417, 5115.8317389664, 
    5084.70344729272, 5033.92500658187, 4967.52780535301, 4795.91350191935, 
    4525.86041312957, 4233.61200905282, 4106.69256570607, 4177.78953786098, 
    4393.32084806382, 4518.35476109077, 4504.83137814346, 4450.12596806817, 
    4399.111723597, 4427.50871686708, 4467.95533467372, 4480.35709656017, 
    4443.35655617591, 4409.05188312619, 4400.65563853428, 4374.27699430758, 
    4375.30473009713, 4381.405747513, 4382.90756996149, 4365.03948381187, 
    4341.0116358294, 4320.29196577935, 4328.40204963706, 4340.51923668607, 
    4332.79164712298, 4321.25855687133, 4343.18398251296, 4349.61767815449, 
    4381.16735337316, 4419.18185522252, 4449.37447965164, 4468.40332626254, 
    4490.28274179915, 4527.36566470826, 4556.77791060894, 4559.72219631862, 
    4509.31747801416, 4447.68359234838, 4362.08607402301, 4278.18572889402, 
    4190.37765881335, 4119.53550763662, 4070.42621396127, 4030.23431148438, 
    3998.3357452112, 3981.46132135912, 3955.97658343563, 3925.08850651842, 
    3878.67766925858, 3817.32412202203, 3761.89754717535, 3721.27612304688, 
    3689.31150249592, 3649.99651825636, 3592.74808984079, 3503.78674192981, 
    3403.79176662216, 3310.68684204702, 3274.50466476914, 3288.54428633844, 
    3298.43442883564, 3276.4970302975, 3223.70969274721, 3189.2289819237, 
    3144.26348834804, 3039.21114266598, 2840.17873838179, 2561.06348997093, 
    2200.83733918469, 1575, 1979.81123140228, 2161.7353516448, 
    2411.66147126736, 2624.06586960288, 2797.28125473179, 2901.53281443914, 
    2902.07602166104, 2758.41088867188, 2558.29366328843, 2272.02244789826, 
    1604.10739395172, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 60, 90, 
    513.14843403502, 1037.63825932765, 1935.05359591651, 2719.38571830012, 
    3356.52979347625, 3767.40844946855, 3992.58154943072, 4116.72137888781, 
    4197.26305134697, 4258.39238392819, 4279.01850753293, 4256.91261520746, 
    4191.16438704538, 4115.36442880452, 4017.32080378702, 3825.41887834037, 
    3680.46835768247, 3562.91195898606, 3540.93105648832, 3595.6653111983, 
    3641.15712983922, 3652.24490937501, 3665.5957549422, 3743.30143480708, 
    3956.68642463787, 4159.84624007918, 4358.57421375797, 4516.79800688168, 
    4615.79738711328, 4622.72510140928, 4528.60121608013, 4399.02420124155, 
    4288.08134708484, 4257.60073200089, 4323.64794547589, 4435.96219294398, 
    4479.40946342898, 4546.23872647494, 4654.49929871957, 4782.61276206324, 
    4896.40342208784, 4966.75126523906, 5014.14111235644, 5053.46335560542, 
    5053.97695865406, 5039.90558504599, 5000.70371633022, 4899.13807784806, 
    4731.83982711223, 4557.79032389304, 4332.99038867443, 4106.49867887069, 
    3750.64603538103, 3345.60795175094, 2776.30284068911, 2327.38623624056, 
    1879.06542324474, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 2515.44003976516, 3159.84831600362, 3632.012385446, 
    4066.34762629395, 4458.81816877942, 4743.55826299292, 4943.31591977202, 
    5029.91779386505, 5033.58797954701, 4960.78453028828, 4824.84384727141, 
    4661.4038787647, 4506.40529941937, 4591.89320915505, 4580.49019669, 
    4548.24233144153, 4462.09963102878, 4331.67009758995, 4156.85700580182, 
    3959.03144636021, 3740.59223531957, 3533.94317367366, 3361.53675224252, 
    3368.65069301571, 3578.76244605589, 3776.18331357237, 3850.3910963356, 
    3593.01857902913, 3052.88711257634, 2640.84402827178, 2989.97012613319, 
    3590.11780735311, 4099.5658266777, 4402.73797726736, 4519.04888974764, 
    4550.33832067955,
  4500.67372456699, 4488.47261213244, 4458.24668699243, 4441.20895026993, 
    4435.70587041734, 4424.94322823397, 4393.30571078261, 4230.75550864506, 
    3967.71248357875, 3643.24995953987, 3749.92468023872, 4091.03924855347, 
    4262.2028378187, 4250.33438615583, 4018.83779355077, 3619.13200395915, 
    3012.03361128566, -0, -0, -0, -0, -0, 0, 40, 40, 40, 50, 50, 50, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 2550, 2550, 2593.35567543021, 2550, 
    2665.35446456005, 2665.35446456005, -0, 1904.35838920445, 
    1904.35838920445, -0, -0, 2268.96343301917, 2692.88965272675, 
    3018.37069488411, 3463.74830367087, 3653.83136494606, 3728.82028992295, 
    3946.4384960009, 4019.28378255034, 4019.28378255034, 4018.68536153038, 
    3837.31074155061, 3556.42785749923, 3346.70275791117, 3371.73008256064, 
    3620.12845499327, 3883.97931271439, 4065.89147763595, 4210.59786396207, 
    4286.93620187412, 4477.02279837461, 4549.62960708528, 4683.80676009411, 
    4574.34318091596, 4173.74994690446, 3622.89089125379, 3074.85053893891, 
    2670.42441141851, 2466.66776221529, 2454.95683012614, 2610.08446453477, 
    2869.3212109161, 3253.803624118, 3686.58945355054, 4039.96644858327, 
    4247.25407332539, 4314.67057251806, 4310.27160566024, 4292.65347679793, 
    4300.35812390919, 4281.42101325179, 4322.40089025465, 4238.19092234936, 
    4174.98439028266, 4053.81920369425, 4118.69210266943, 4399.01684284677, 
    4688.85979555522, 5035.07386468381, 5284.55991066076, 5395.1735236335, 
    5413.19637120084, 5329.01221745204, 5296.64734627135, 5241.4436966787, 
    5212.10853704358, 5295.58683913812, 5358.17074536295, 5436.97016743764, 
    5451.76816170284, 5444.22238019551, 5435.49193406395, 5405.32309925541, 
    5354.66241924743, 5305.81258133785, 5260.38398283592, 5205.30706131609, 
    5150.30746108908, 5090.74626883308, 5023.85758260173, 4936.48898383907, 
    4725.30800664573, 4421.10934467257, 4129.14858842125, 3972.05404809528, 
    4146.01910097422, 4399.13417725031, 4521.86051709788, 4516.94677794981, 
    4471.79830400336, 4426.36936466239, 4453.79106585846, 4501.22930190158, 
    4520.19022075177, 4481.57696792021, 4445.11024662749, 4424.84922093479, 
    4391.91070069528, 4388.43426920216, 4385.30473971934, 4387.91710292287, 
    4369.79309595398, 4341.73000902586, 4321.65310880571, 4327.66825713453, 
    4343.17605967145, 4346.81344011636, 4339.36323581749, 4347.70594221237, 
    4346.32730812943, 4379.61161628635, 4419.34957546162, 4448.8901757492, 
    4466.51056380692, 4485.35162896448, 4521.99189862539, 4558.65822778385, 
    4567.07499168683, 4519.55598532965, 4460.49189120846, 4373.94035642779, 
    4291.36137796471, 4205.33289976948, 4126.81829644149, 4065.89147763595, 
    4018.17239887886, 3980.46697092547, 3961.3497916675, 3932.86774698744, 
    3905.18329521175, 3864.1232061479, 3809.38778527081, 3758.37529968078, 
    3721.27612304688, 3687.39115206496, 3645.3722604175, 3585.75954364839, 
    3500.04580608866, 3400.74817706678, 3310.42809935428, 3273.22812645036, 
    3288.74830732632, 3295.66684640582, 3267.35659797965, 3201.26859625955, 
    3160.75928891502, 3101.95758218984, 2987.07994969387, 2804.79058919041, 
    2519.35703643531, 2219.12659563441, 1650, 2011.7722151717, 
    2201.3540617624, 2434.85843211172, 2645.54881692062, 2826.69519478631, 
    2943.96572199995, 2955.27304467894, 2824.19962568481, 2638.42343361752, 
    2357.23100199984, 1657.07516731982, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 80, 170, 629.3616004902, 1289.0608245216, 2225.79923667399, 
    2963.55521086378, 3522.62657548162, 3898.54848611874, 4094.42043673199, 
    4184.26636641796, 4244.72625239133, 4261.30906260115, 4276.26055813709, 
    4236.72076238626, 4148.49922924405, 4045.07256738348, 3916.30637890694, 
    3721.27612304688, 3567.41690836512, 3450.23684911743, 3472.71911741798, 
    3549.47712392797, 3639.20368873357, 3656.98767499962, 3695.71311984587, 
    3769.01611130578, 3992.15929096539, 4202.24970742118, 4385.71685300404, 
    4543.21513212247, 4655.33124939481, 4688.19534506528, 4645.63000022703, 
    4535.39210379056, 4429.35933086565, 4365.94745515626, 4419.18185522252, 
    4500.26885652522, 4534.03081211137, 4589.05278819452, 4675.20328891006, 
    4779.07571895829, 4859.45211892486, 4934.41665178681, 4980.24007372586, 
    5012.23590377359, 5016.15009456976, 4989.56024515303, 4967.44115577564, 
    4895.22691545502, 4725.37695201388, 4548.49860307981, 4324.54636383105, 
    4085.73648841755, 3702.83488875433, 3275.7236660768, 2758.41088867188, 
    2218.5094383242, 1838.76493502209, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 2296.72918486572, 2961.68545488931, 
    3479.54834932689, 3966.75791317459, 4336.65074504388, 4669.89009468053, 
    4905.91508255781, 5023.00565395588, 5044.95372457558, 4978.00004697137, 
    4857.58574159541, 4712.73522775228, 4550.25053521458, 4593.61975158299, 
    4572.98134954829, 4530.2589028152, 4435.32491260525, 4287.72878100702, 
    4094.96705092812, 3894.57261692134, 3665.1588948581, 3484.32312429983, 
    3333.27237766794, 3376.59782254459, 3606.24637209221, 3807.00532059276, 
    3859.34350030905, 3557.297640502, 3012.04483329963, 2600.59225354976, 
    2876.25854540909, 3469.09285599527, 3997.90364869059, 4310.29740561477, 
    4446.19282430846, 4486.51434604212,
  4461.47037414104, 4450.36941410168, 4426.86635621506, 4419.18185522252, 
    4401.33116349405, 4385.21477344037, 4359.2848459265, 4213.29922001113, 
    3941.34606497926, 3524.53992009984, 3571.76658946419, 4107.41415347489, 
    4192.88179221167, 4146.76280882106, 3910.74299447357, 3622.83289689466, 
    2718.95316328772, 1136.76173782374, -0, -0, -0, -0, -0, -0, 40, 50, 50, 
    50, 50, -0, -0, -0, -0, -0, -0, -0, -0, -0, 3300, 3300, 3300, 
    2966.47399291501, 3290.64660247986, 3237.21752635682, 985, 
    1891.04361589842, 1891.04361589842, 0, -0, 2846.585140864, 
    3077.71160570778, 3290.69446831092, 3597.44647894483, 3787.73243388295, 
    3861.76623364374, 4073.85712360613, 4153.28605769625, 4230.43625088683, 
    4168.92373306701, 3934.74231067321, 3590.27143207269, 3281.82806417706, 
    3354.22817653202, 3745.07378228933, 4054.1793933575, 4237.52071694129, 
    4339.50381380426, 4373.41898472792, 4670.54344167102, 4589.20652033612, 
    4595.25764708187, 4619.34065417279, 4152.06193306475, 3632.42137162029, 
    3086.1207068686, 2702.8612853673, 2519.46291859642, 2523.30460120844, 
    2682.1022488691, 2893.50122543634, 3289.52726262524, 3721.27612304688, 
    4065.89147763595, 4259.06627536323, 4304.58239204041, 4299.87852886115, 
    4291.86147206055, 4323.62386537217, 4270.64649533259, 4344.84831495176, 
    4242.40327379544, 4189.98378957422, 4028.85314487633, 4065.89147763595, 
    4399.01684284677, 4753.39579071224, 5043.84332923614, 5324.67838464455, 
    5416.78679295781, 5429.35421847326, 5388.77481496634, 5305.90519687777, 
    5170.83158724948, 5264.2730095512, 5307.01131285244, 5374.52145374104, 
    5440.24831023059, 5441.90152962071, 5426.89673301032, 5440.29415500638, 
    5389.14167890948, 5354.58967628343, 5332.66607409202, 5294.48723432025, 
    5227.55502117396, 5175.26496234147, 5115.37959329741, 5037.66911876662, 
    4940.01271470195, 4723.9191917212, 4335.52432296548, 3996.562263644, 
    3621.53181203824, 4121.11630421913, 4450.47597482384, 4537.33528490203, 
    4564.36139186165, 4480.56223576169, 4419.54010627078, 4470.42042351422, 
    4562.34146531537, 4573.4852817499, 4519.73658145478, 4489.84863377964, 
    4463.08264532313, 4404.90426702358, 4397.76588461657, 4389.34378959349, 
    4393.27022449429, 4378.30897569649, 4334.97663634171, 4322.49414940367, 
    4326.03620639198, 4356.35369974203, 4377.59262765165, 4366.48887952371, 
    4366.14381884484, 4331.44401155524, 4370.53526953382, 4419.18185522252, 
    4449.65933236906, 4472.3820374204, 4468.67730456425, 4508.97693505483, 
    4570.33555372926, 4590.89191155707, 4535.88507271322, 4483.55806017677, 
    4387.22487103913, 4324.16422141219, 4238.02652923784, 4139.46819903543, 
    4055.69324190393, 3998.78502738653, 3953.79276854743, 3939.11274627238, 
    3898.4647503186, 3886.37618485382, 3845.01066233681, 3799.38720865469, 
    3750.98498214615, 3705.39307198126, 3689.83809861644, 3639.18170925316, 
    3573.62506934696, 3496.17922988966, 3395.9771047528, 3298.63472407642, 
    3245.05209241594, 3295.36785360755, 3300.84643887038, 3266.30272783858, 
    3153.15221044076, 3133.50399658274, 3049.98990832176, 2928.15245630122, 
    2758.41088867188, 2494.456372955, 2230.59305265195, 1785, 
    2096.04474509645, 2280.66705127646, 2477.89220397105, 2663.08670316444, 
    2814.69283326296, 3003.73541314293, 3003.73541314293, 2930.9666361283, 
    2772.75091036104, 2531.33418932142, 1657.07516731982, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 110, 307.862556489688, 686.627904008391, 
    1554.16343620012, 2588.27842026556, 3310.45448686455, 3756.0699438644, 
    4065.89147763595, 4175.31170693102, 4260.26985849912, 4280.87036421438, 
    4233.85998030403, 4272.37563942844, 4184.8659737215, 4119.10434175367, 
    3958.77930455623, 3796.59386619614, 3577.28642127358, 3432.70762591016, 
    3290.5456338665, 3421.48301899893, 3495.91474781455, 3643.17534306633, 
    3650.12914137371, 3729.86908422183, 3728.77141233092, 4065.89147763595, 
    4256.86804838188, 4443.02177718588, 4578.7836179576, 4715.21993248963, 
    4740.23614604055, 4740.23614604055, 4695.07306093343, 4656.33216980602, 
    4496.89475451454, 4557.73200936542, 4577.41698489989, 4599.13462913121, 
    4671.80987327315, 4708.63040913516, 4698.61309389974, 4813.30794650173, 
    4885.10618111404, 4938.18246501891, 4967.3280206481, 4944.43200303872, 
    4969.64230040766, 4949.09289515972, 4865.0527931547, 4713.03454514226, 
    4549.40237256381, 4326.72760623346, 4065.89147763595, 3640.31595004329, 
    3229.55606009627, 2732.67662831083, 1940.6265026171, 1872.22652234516, 
    994.228752204076, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 1629.24516766314, 2626.68260308271, 3314.9764301273, 
    3858.17488621377, 4247.76988295988, 4580.26698918709, 4890.21202621084, 
    5014.37940013758, 5061.94357993825, 5018.92082127192, 4904.30690921522, 
    4779.07571895829, 4595.98509987755, 4597.57105754736, 4554.83085929122, 
    4515.14811964854, 4419.18185522252, 4226.31790353223, 4033.75745271511, 
    3825.09537406128, 3591.98969718421, 3428.56626510957, 3264.15248551606, 
    3376.59782254459, 3660.83926561322, 3871.58552319473, 3888.45535845882, 
    3592.03474474194, 2978.38797919796, 2466.66776221529, 2700.41072427266, 
    3333.60682136821, 3897.4726594857, 4242.2004146105, 4370.61631687186, 
    4423.37836666829,
  4419.18185522252, 4419.18185522252, 4391.92045176035, 4377.28356002389, 
    4360.10686948764, 4340.96496907364, 4304.34804454936, 4164.00375808304, 
    3847.29618354355, 3413.68761240594, 3505.0495456418, 3976.29832953288, 
    4032.89580106251, 4032.89580106251, 3776.53354418548, 3338.91600390563, 
    2081.15247247426, 1136.76173782374, -0, -0, -0, -0, -0, -0, 40, 50, 50, 
    50, 50, -0, -0, -0, -0, -0, -0, -0, -0, -0, 3300, 3575, 3587.85201512091, 
    3749.23260314192, 3970.76958225497, 3952.57445416344, 3205.32548130156, 
    1891.04361589842, 1905.71712968336, 1905.71712968336, 0, 
    3125.87240225461, 3453.21067924662, 3645.58088493152, 3587.87949574083, 
    3857.87258045954, 3946.52627371475, 4184.82709587917, 4269.22776755674, 
    4323.8415465999, 4227.6428114055, 4005.35662813926, 3657.49551869394, 
    3247.99334744559, 3408.18957701359, 3859.92538010013, 4151.9670354406, 
    4343.42531148712, 4419.18185522252, 4446.18094319598, 4711.65216869178, 
    4595.84411891614, 4766.42491482815, 4595.25764708187, 4168.92566090139, 
    3641.01907911815, 3096.61690362743, 2760.14430551101, 2590.75779093039, 
    2635.32795405865, 2758.41088867188, 2968.11058005494, 3329.61391730534, 
    3721.27612304688, 4065.89147763595, 4258.11293120709, 4298.67512092404, 
    4294.36219943157, 4287.27127174526, 4334.47934523396, 4286.42121628379, 
    4323.79142085279, 4188.06818681973, 4163.5013117641, 3979.42691184733, 
    4046.65637028433, 4319.9052743737, 4827.98228604807, 5070.30727292577, 
    5340.4954341412, 5425.63844769253, 5450.47096731979, 5395.58061151684, 
    5327.86404327077, 5261.89043065856, 5263.84972845676, 5240.26682541121, 
    5355.33462486798, 5447.06394147121, 5427.88066741815, 5407.67103321436, 
    5411.29243654436, 5374.01213146067, 5382.65904365707, 5345.50319760866, 
    5326.14459112234, 5241.21403963204, 5026.38657730104, 5110.23355060996, 
    4959.46299642966, 4857.48656990748, 4606.69445351343, 4250.09966154897, 
    3844.87198893088, 3409.70955175411, 4145.12779051088, 4502.37233355872, 
    4606.51350844776, 4641.58726294458, 4561.19763267473, 4513.39815066852, 
    4541.8889114465, 4632.2622575572, 4644.71954501715, 4588.52081032366, 
    4549.42751725101, 4492.4539226536, 4439.36411972752, 4422.26035708647, 
    4397.18403940978, 4407.01730052175, 4380.01420929001, 4340.09447322869, 
    4308.01218506614, 4333.47686684824, 4345.02300004776, 4369.43989562816, 
    4361.62281064735, 4372.73288785875, 4348.94933191097, 4384.15494174847, 
    4419.18185522252, 4436.24879014232, 4462.60762445727, 4462.51457968966, 
    4522.32702796438, 4556.51145389999, 4586.6421559514, 4545.75554353315, 
    4489.3864092514, 4396.70627869742, 4316.70146240958, 4251.31526708949, 
    4158.21113889544, 4086.2287114533, 4017.26174276577, 3965.14101088221, 
    3921.60834257087, 3879.00374383542, 3865.51649288811, 3832.54773965999, 
    3798.61227990743, 3761.82951974735, 3735.86017978729, 3698.945798199, 
    3642.77382699203, 3569.2011928851, 3500.69646827401, 3401.05284500429, 
    3285.88516489882, 3299.56269795911, 3240.68761047056, 3213.89847893116, 
    3179.92897604663, 3091.55355856045, 3044.86391559682, 2966.59799981692, 
    2864.14546918625, 2708.7255482979, 2481.92528863878, 2274.9367200949, 
    2120.13474438469, 1919, 2318.84397117162, 2475.4036921477, 
    2675.79594120517, 2818.29714087672, 3013.6032315099, 3004.86195345535, 
    2942.20184014914, 2783.69634203585, 2559.08561659346, 1871.7611272836, 
    1115.34121330582, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 60, 110, 
    393.228739433858, 858.239647084743, 2005.67458759425, 2902.97936094534, 
    3524.23188513666, 3929.24236766206, 4149.37100096462, 4234.70669817089, 
    4300.53773369352, 4330.16178733568, 4337.43616427442, 4289.51924343266, 
    4172.02407358469, 4105.95223102656, 3940.14778974323, 3721.27612304688, 
    3500.84423840564, 3307.901832865, 3209.35431482732, 3411.88036874402, 
    3510.68554988855, 3668.07554207837, 3755.83838167586, 3850.93635390197, 
    3846.46631156421, 4096.64125159182, 4239.94033385745, 4443.59840271962, 
    4591.06895385108, 4715.21993248963, 4837.59942914786, 4825.65989744821, 
    4794.46026919174, 4760.27320087605, 4602.68649541612, 4655.31097002499, 
    4625.2649771758, 4557.9225139907, 4571.86064118803, 4593.65732640997, 
    4686.27312199962, 4646.8921322852, 4746.37692614592, 4805.44464576777, 
    4830.43450299381, 4825.23212252256, 4826.9001464491, 4849.08576869787, 
    4809.73079923265, 4685.29655254082, 4509.92418215603, 4294.68786049152, 
    3989.40098897418, 3552.70995225529, 3106.68871581075, 2656.12058969289, 
    2134.86900396266, 1858.63937124456, 1170.70609572657, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 1961.97468079322, 
    3038.02832469574, 3619.42962499743, 4077.00445800893, 4441.08214963292, 
    4822.88830309258, 4999.46660893168, 5058.51540536626, 5037.10721423967, 
    4941.65911708396, 4840.06557371929, 4680.84004242418, 4606.52877572644, 
    4571.56085720396, 4514.68479200253, 4356.46929896766, 4186.71106452269, 
    3912.02146619238, 3776.7985513156, 3545.11361631838, 3350.08686994658, 
    3218.47209626472, 3450.25431121424, 3706.05974323447, 3880.08888596237, 
    3897.70008875766, 3567.80062200883, 2927.78423161869, 2163.65344429691, 
    2607.87582267341, 3221.0951180781, 3788.76109287423, 4130.49084476188, 
    4201.08267832746, 4357.92275363666,
  4357.38273788739, 4381.03465004424, 4361.50944703394, 4335.95700226493, 
    4315.71498761982, 4293.90691721381, 4235.94663010972, 4107.70076828297, 
    3822.04143468451, 3484.40801911152, 3463.81645218572, 3849.6095106815, 
    3945.77315957503, 3824.77308386006, 3396.7543394752, 2627.17713375318, 
    1850.02248997134, 1151.61501345749, -0, -0, -0, -0, -0, -0, 50, 50, 50, 
    60, 60, 60, 60, 60, -0, -0, -0, -0, -0, -0, 3300, 3575, 3747.56921169544, 
    4171.59026742216, 4281.91522360047, 3993.63642988682, 3339.9012273508, 
    1520, 2143.85575351396, 2307.24928560866, 2449.33311410393, 
    3172.76862012086, 3535.59228801862, 3641.75754405651, 3742.11539634606, 
    3905.64274313015, 4084.18734470563, 4264.57345654197, 4361.99436024138, 
    4386.51763778297, 4239.21422325664, 3996.52890504007, 3668.9024094139, 
    3332.7907027525, 3436.67263372042, 3808.03670914984, 4135.66349675512, 
    4341.53333884411, 4421.42978772972, 4463.12222367644, 4588.10760264682, 
    4611.75183996093, 4710.41846629413, 4536.31909034967, 4154.20868986485, 
    3683.62151779159, 3176.6909244118, 2863.86450281457, 2723.21101904309, 
    2748.13823347331, 2870.26545479895, 3065.78548661781, 3411.32316264811, 
    3739.51881126413, 4036.31162215805, 4239.53698703814, 4304.43973166023, 
    4326.74149346836, 4333.95061333416, 4350.86594949929, 4328.7919528259, 
    4296.95975878654, 4193.45857949493, 4133.83119298121, 4075.41997403038, 
    4178.19936104953, 4456.85548802496, 4836.41446567181, 5125.24317239387, 
    5352.34315366582, 5441.01536770496, 5458.48780126217, 5403.81234497126, 
    5333.45376917159, 5265.00680299484, 5237.75939899514, 5226.92467933201, 
    5298.70023089871, 5379.559721852, 5391.9351331107, 5412.48418685488, 
    5418.31865349341, 5408.00395237689, 5385.47765627905, 5363.16635052421, 
    5320.0996786452, 5230.57284805417, 5130.76260297652, 5070.99193032119, 
    4942.98605446463, 4745.54285964629, 4441.31325986937, 4065.89147763595, 
    3751.62819983205, 3854.4533677897, 4211.36576926922, 4500.35605485138, 
    4641.49118777882, 4672.46194033115, 4641.34370325581, 4622.97418444704, 
    4632.67924154743, 4682.93321966714, 4690.98998665337, 4650.45425046203, 
    4599.6538144985, 4547.39364627638, 4489.12938269885, 4457.29474919143, 
    4432.76867157623, 4419.18185522252, 4377.31860702514, 4348.4341147669, 
    4324.29304759784, 4339.7652664777, 4348.84387720572, 4363.93810776499, 
    4345.96566380166, 4365.01750677946, 4359.75086810608, 4383.12002591573, 
    4419.18185522252, 4442.4576962777, 4458.08494684715, 4466.70964743568, 
    4506.31013550694, 4536.80293313767, 4546.4185297058, 4518.95181399788, 
    4464.73436496913, 4394.28171712686, 4311.03873527864, 4237.08562865696, 
    4170.65848451071, 4101.98077987403, 4036.95071207797, 3978.58900929569, 
    3922.25552394315, 3885.14311590637, 3870.30919583259, 3838.52698206735, 
    3808.83240449258, 3780.85040716835, 3750.2995136216, 3721.27612304688, 
    3652.50269989286, 3579.09481136449, 3502.83764475735, 3398.89789112674, 
    3306.98183820233, 3284.31639836014, 3258.29626867629, 3239.1053966654, 
    3189.0467844081, 3139.52233197032, 3092.51004380698, 2996.41698588494, 
    2882.78931046649, 2747.36161807917, 2572.59088685163, 2397.20103137894, 
    2246.82038838901, 2191.85384798669, 2261.72919112702, 2433.24949484485, 
    2625.99047537464, 2828.4219358319, 3004.86195345535, 3004.86195345535, 
    2902.42511457794, 2758.41088867188, 2567.37192247777, 2260.8311087775, 
    1511.15189479409, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 130, 294.462890625, 
    596.260553944861, 1205.09233171499, 2213.88155215359, 3027.95991220103, 
    3623.64958000038, 3984.65253499972, 4177.97462345693, 4249.50344127261, 
    4298.93716651105, 4348.35792192317, 4343.59196379839, 4280.65332261218, 
    4159.46531153025, 4040.436968937, 3873.53568172009, 3657.86748722896, 
    3437.58202480956, 3281.18423924381, 3264.04490223828, 3419.52949624078, 
    3562.57311333671, 3723.24999383541, 3838.20064678319, 3934.35508680016, 
    4002.92873509327, 4142.58068692625, 4259.47038603371, 4387.89780719885, 
    4528.69213078143, 4709.99961381393, 4842.10274659261, 4859.68099022066, 
    4819.0687079493, 4762.84490677225, 4657.91461289738, 4650.0669680746, 
    4601.81570555949, 4550.10000896927, 4478.29484125613, 4425.84123949975, 
    4508.31558103849, 4524.55197325715, 4548.50691784466, 4578.85978442575, 
    4564.4271109357, 4590.59029744464, 4610.77964816295, 4644.71304689528, 
    4597.15106405018, 4560.94458378024, 4424.80056146343, 4187.86953656124, 
    3842.16925837656, 3363.42459158802, 2873.41954194069, 2407.06976664592, 
    2002.73252841093, 1708.37172826823, 1184.62222704214, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 2701.80846770991, 
    3347.95817436827, 3839.7912368812, 4272.08238116926, 4703.96864157866, 
    4938.11989119244, 5035.09798859796, 5028.19545400166, 4935.21936434778, 
    4846.6174870216, 4704.07353849479, 4596.72112803616, 4554.71230131454, 
    4471.06264934651, 4298.89344927439, 4083.37753806057, 3831.34594798656, 
    3661.58907774832, 3443.44268331537, 3301.9696553252, 3277.19483767084, 
    3470.3321121232, 3721.27612304688, 3882.819446979, 3863.44327723064, 
    3477.29199130538, 2849.53708187536, 2323.53236020221, 2576.70455623396, 
    3095.40997025206, 3649.09055794278, 3959.05932938739, 4071.64754201871, 
    4273.24435315215,
  4301.93617353715, 4340.85471279668, 4325.40215661622, 4295.21381111623, 
    4271.76660167632, 4249.71679781118, 4198.58132977571, 4068.29729406405, 
    3796.98719033241, 3474.75266041418, 3417.94372611667, 3750.0419290348, 
    3809.35057806939, 3596.68103296748, 2988.06489195354, 2230.67840315254, 
    1605.45970138867, -0, -0, -0, -0, -0, -0, 0, 50, 50, 60, 60, 60, 60, 70, 
    70, 70, -0, -0, -0, -0, 0, 3300, 3575, 3831.0587220944, 4348.98352268653, 
    4330.75758910167, 4165.66114142338, 3498.10025046266, 1450, 
    2348.54384633699, 2560.62168282655, 2900.90236576543, 3474.23489745566, 
    3725.07832936719, 3751.94626411642, 3793.50841464248, 3962.7565340701, 
    4148.65649928903, 4320.25952355233, 4403.36582580491, 4403.36582580491, 
    4281.33615433514, 4032.70718179633, 3695.75068189956, 3353.62078527875, 
    3433.47841849433, 3799.3559749153, 4137.5650435056, 4337.28784423564, 
    4401.65224956243, 4435.66088543911, 4498.33089273407, 4570.75244123011, 
    4673.61999852747, 4517.60882319307, 4159.34554211427, 3690.55659763628, 
    3237.37730939095, 2947.9259287168, 2822.79589639755, 2850.3090848137, 
    2973.92636596661, 3179.52584967316, 3483.17934501814, 3765.30188675433, 
    4040.45806274117, 4239.52092053726, 4323.45195324797, 4361.3086151944, 
    4372.19670985122, 4374.05339890388, 4336.32876567271, 4294.66807191186, 
    4197.6747825806, 4137.51848706566, 4072.59475431192, 4250.57192633453, 
    4546.14091090844, 4888.26382771879, 5157.42757736263, 5382.33527344328, 
    5463.33674277186, 5485.26136622647, 5434.05304182655, 5343.4828615311, 
    5262.95530878301, 5216.05751394257, 5212.35575421184, 5273.6692208731, 
    5332.45794140689, 5385.18347303105, 5412.27644493148, 5429.25369643427, 
    5432.62178826406, 5388.23189763356, 5369.72109588198, 5328.51578284321, 
    5222.81696023481, 5126.08012352739, 5029.28467573826, 4862.47683194122, 
    4603.92049127819, 4302.81043301608, 3935.96868842057, 3698.16294464861, 
    3950.80317510031, 4253.22925866367, 4522.79028284897, 4682.34524116754, 
    4715.14810564224, 4708.97433802882, 4712.93673582068, 4729.94285912427, 
    4757.87783937146, 4750.08580976035, 4710.20829563428, 4658.09067831441, 
    4601.07627477804, 4539.13582856955, 4493.16957781751, 4461.19750832982, 
    4426.06034302654, 4385.62744893972, 4358.25426764117, 4338.000998397, 
    4354.02817653389, 4365.31980779237, 4376.91336878568, 4354.2951020201, 
    4372.60729426346, 4365.10409815315, 4382.77588362316, 4419.18185522252, 
    4438.9003086047, 4451.61488121468, 4461.8315108834, 4494.19283656416, 
    4517.84223804007, 4526.53884740281, 4503.20878924633, 4449.11035345648, 
    4380.70126945464, 4308.10624590163, 4236.33714188289, 4178.95266887203, 
    4118.05114753243, 4065.89147763595, 3991.92473455131, 3928.59504278483, 
    3892.5341652581, 3876.86699670806, 3852.84501332496, 3827.72684452454, 
    3800.01902886831, 3768.82522977269, 3729.95923369335, 3667.59885058037, 
    3592.0032723691, 3504.44309769543, 3399.55669263503, 3306.50815151161, 
    3283.43594561796, 3277.56066382934, 3270.54102310698, 3228.22770893511, 
    3203.45441121861, 3155.64666602018, 3045.82527459837, 2932.81775849485, 
    2804.34106517033, 2663.54907686761, 2492.73442563659, 2339.47225876876, 
    2238.3522861058, 2218.95472845005, 2357.48729633917, 2560.20041149779, 
    2787.53943464943, 2968.14864888051, 3025.87941648547, 2882.49571987416, 
    2758.41088867188, 2594.39435095417, 2410.91983706194, 1757.86190739015, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 140, 454.636363652683, 
    803.625015916513, 1482.71199164271, 2445.81226181486, 3208.93690930273, 
    3751.72194186795, 4067.92091552841, 4199.721162969, 4263.72076968913, 
    4306.45461178203, 4362.38137340341, 4355.9308323953, 4275.85080171382, 
    4147.70269034774, 3997.03532512898, 3806.25774387936, 3588.99142579313, 
    3376.79951834829, 3237.18721042602, 3277.68577597718, 3449.99393868464, 
    3615.71220542939, 3793.38741775636, 3925.25938663608, 4030.53436115963, 
    4096.80853754669, 4189.24610759061, 4236.23744056007, 4338.69624771872, 
    4468.2051835596, 4672.03310044817, 4845.43374218072, 4882.06409508149, 
    4853.82273058852, 4804.67283934928, 4719.39497712977, 4655.36284174476, 
    4557.80514562072, 4460.49714471375, 4308.8494046354, 4276.65903710714, 
    4287.64625626269, 4344.97605568358, 4345.27259251888, 4347.47144220056, 
    4301.09061834633, 4350.8507065856, 4405.8920006908, 4474.7391695763, 
    4434.1991527653, 4391.15156325741, 4318.30066946376, 4065.89147763595, 
    3655.91952804144, 3177.69961734332, 2629.58541241101, 2143.40291412915, 
    1818.65709506208, 1542.03948663489, 1184.62222704214, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 2388.03779399053, 
    3107.3156703982, 3633.81290910997, 4099.89074674153, 4573.81678118793, 
    4883.91042922426, 5016.6546668292, 5029.9188992603, 4952.80130984023, 
    4864.27086704334, 4731.42137308214, 4600.44698189626, 4523.10000389368, 
    4419.18185522252, 4202.81485794346, 3978.09211278708, 3736.01160924375, 
    3568.63902963492, 3392.96671856764, 3306.11568018447, 3307.4440877051, 
    3498.0255712046, 3733.99455401208, 3903.93728825089, 3845.36657270762, 
    3441.90873070594, 2758.41088867188, 2222.78645735042, 2516.30672226209, 
    2975.38732573928, 3518.40312990781, 3802.29075151395, 3962.33115382049, 
    4194.85757630828,
  4244.13210224914, 4290.79411304315, 4287.71969717677, 4257.81837670703, 
    4231.68238149382, 4209.20553017545, 4167.25104412612, 4039.63625064965, 
    3787.88888927184, 3480.97213824518, 3387.2978515625, 3681.22971735439, 
    3709.71615838002, 3394.03440289519, 2619.06754861085, 1944.05364782763, 
    1450.5465508743, -0, -0, -0, -0, -0, -0, 0, 50, 60, 60, 60, 70, 70, 90, 
    110, 110, -0, -0, -0, -0, 0, 2359.85387208075, 3246.14735692727, 
    3825.63250567852, 4330.75758910167, 4330.75758910167, 4273.31290072133, 
    3619.68847873104, 1450, 2348.54384633699, 2758.41088867188, 
    3283.52248773559, 3789.15321139376, 3901.70938794606, 3861.84574379022, 
    3850.39384446278, 3974.76385591515, 4217.59581182274, 4383.22091571693, 
    4456.6955223597, 4439.50604178342, 4310.89596431383, 4073.10084182052, 
    3722.86224660104, 3341.62609234643, 3416.36424653216, 3775.3014416549, 
    4114.61447095533, 4319.00251617269, 4371.02672092098, 4377.2859556821, 
    4419.35170919185, 4532.79232137588, 4610.14405900841, 4476.01134213311, 
    4151.5770009682, 3721.55268768493, 3279.92950536544, 3021.25300320536, 
    2913.36050769864, 2929.64364250758, 3068.23796431694, 3294.80829818021, 
    3548.24686564841, 3782.89474132991, 4054.59156538795, 4260.59607938885, 
    4350.44738921693, 4407.7245321105, 4407.7245321105, 4402.40660408906, 
    4344.28019023002, 4274.66200522438, 4204.30911713627, 4145.83748064151, 
    4091.35743501526, 4304.37229668287, 4631.87280772618, 4942.44090523994, 
    5189.45888581798, 5414.32620729858, 5496.70912042421, 5500, 
    5460.45809255079, 5353.28414179956, 5265.18566695815, 5185.29910328721, 
    5189.85624621291, 5259.44036544058, 5315.58328752256, 5381.56113294134, 
    5419.15191494155, 5446.45164999886, 5460.34827849467, 5400.27341124148, 
    5373.48925606834, 5322.14337950556, 5224.0456812312, 5110.7795111467, 
    4976.13168111781, 4743.40910425308, 4473.04810960197, 4166.24742212751, 
    3809.15386244751, 3710.74266912742, 4025.98653661611, 4300.07461713566, 
    4544.47800648817, 4698.64110666497, 4746.36513866543, 4756.76498964535, 
    4783.68527551256, 4808.35564152049, 4826.26167692363, 4807.12992277879, 
    4779.07571895829, 4713.13000488903, 4654.92068696035, 4587.51718236622, 
    4524.64459007451, 4484.83388176726, 4444.16974224648, 4398.11523783678, 
    4370.242008974, 4355.63780862762, 4373.89025415788, 4384.25935819075, 
    4387.54008411648, 4367.2348235056, 4378.55366790719, 4366.0915395627, 
    4383.51615180171, 4408.16392555798, 4431.31251171723, 4443.40165393816, 
    4457.66348774287, 4483.55580939567, 4497.92319704629, 4507.29869248172, 
    4486.08085287427, 4434.60110861436, 4360.69159057539, 4299.11034883072, 
    4234.36727438841, 4186.04681311506, 4132.71302125383, 4077.58592501925, 
    4008.73252734186, 3942.12488832819, 3904.76735609389, 3889.15341668545, 
    3871.10837639243, 3847.9878091621, 3818.23330595019, 3786.07153011158, 
    3747.65493857407, 3685.57678370652, 3605.96420430466, 3502.08595882728, 
    3398.37872338126, 3300.74742695077, 3281.40548686937, 3293.51838518161, 
    3302.35608892193, 3280.67711161271, 3270.48415351744, 3222.40558860269, 
    3115.66418100574, 3004.1401359601, 2887.13604088013, 2758.41088867188, 
    2606.70543619572, 2436.19862091155, 1785, 2201.15992184028, 
    2274.69253518629, 2479.36351269377, 2742.85400852008, 2933.33276908236, 
    2990.40628588641, 2862.64665033316, 2712.58387997662, 2595.54348007828, 
    2513.82449532961, 1996.33690394119, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    140, 612.432103402777, 1019.71415885479, 1741.82131617511, 
    2643.4515198774, 3337.62835714341, 3847.5663348448, 4087.94952612712, 
    4191.35744053944, 4239.21130546382, 4306.03483424871, 4376.68078780146, 
    4369.84565953189, 4282.11312423237, 4145.62567825318, 3972.76925594098, 
    3756.25294330922, 3532.85514196345, 3334.6883118688, 3216.0064321398, 
    3312.33614265873, 3502.41524998613, 3677.79696773154, 3862.29727700319, 
    4000.43630757956, 4105.27588011736, 4171.8543803232, 4208.28922255151, 
    4185.83526679204, 4251.06521710388, 4389.63561253473, 4621.58294470194, 
    4830.16763066955, 4904.67812615477, 4892.52816189714, 4834.69584710171, 
    4754.88215156913, 4650.85920009511, 4513.09924045916, 4331.69044599359, 
    4169.70853145877, 4096.14001592353, 4049.33958931032, 4088.25415802981, 
    4134.88455291127, 4128.87714819655, 4100.97313791271, 4084.75063064774, 
    4102.33087259449, 4215.43869408002, 4231.49415781462, 4168.09170150351, 
    4098.24369255877, 3859.25387162932, 3489.15433229475, 2976.02438014049, 
    2353.49792766815, 1847.26308919629, 1593.50175536015, 1305.72529879764, 
    1023.9902654882, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 2244.88479703199, 2826.43331408494, 3420.83689089622, 
    3934.9285889491, 4460.71197426439, 4841.27819914199, 4997.66435400116, 
    5027.91943232524, 4964.30483573383, 4865.25088342513, 4729.40389579077, 
    4604.57974529996, 4487.1634722171, 4353.43490228766, 4115.00984070949, 
    3882.52587167371, 3641.80674812859, 3486.99693580825, 3387.2978515625, 
    3341.20831481447, 3372.77702807811, 3543.71686099423, 3762.33737762097, 
    3921.07994592571, 3830.04419508895, 3413.74505232204, 2685.62078684018, 
    2131.55069829809, 2466.66776221529, 2884.86527958765, 3393.58633321442, 
    3662.62091920846, 3864.38292467866, 4130.5907048841,
  4122.27651474962, 4185.01241316976, 4206.46536310333, 4212.6910735063, 
    4180.60410767831, 4155.75577675078, 4126.82987183979, 4007.21356165157, 
    3771.03341617247, 3473.75601585417, 3353.82763717925, 3591.81887352044, 
    3579.12191082704, 3108.17852851653, 2331.946878309, 1744.34306108543, 
    1222.13659397283, -0, -0, 50, 50, -0, -0, 50, 60, 60, 70, 70, 70, 100, 
    130, 180, 180, -0, -0, -0, -0, -0, 2135.99638987546, 3040.83426627928, 
    3672.42683702324, 4241.39383042, 4337.40789742607, 4337.40789742607, 
    3787.48574735902, 1766, 985, 2924.06037155598, 3688.32324180599, 
    4119.05809503975, 4123.72799700884, 4028.0697099851, 3907.04361222971, 
    3977.56275204079, 4272.49290098818, 4466.11712029552, 4510.78108483832, 
    4469.91025243957, 4336.10090042898, 4104.85317959806, 3746.6183876405, 
    3323.6332938013, 3374.46733946682, 3721.27612304688, 4054.90761577172, 
    4269.06247583793, 4303.18848764822, 4282.97939277241, 4297.03041698937, 
    4443.03070057622, 4495.69986825374, 4399.91696917581, 4156.54140498377, 
    3760.28193929925, 3358.29750997081, 3136.17709936001, 3053.59926402898, 
    3028.98827017531, 3170.78521741086, 3426.52476465233, 3633.18273967286, 
    3824.22619269459, 4095.89135082939, 4303.98122570574, 4419.18185522252, 
    4478.4446512194, 4472.66862409551, 4444.08296761405, 4329.67539962061, 
    4267.72665605821, 4185.44198283656, 4164.13556148175, 4118.69113296096, 
    4379.27694640822, 4716.63469204842, 5002.45071304067, 5243.67464250429, 
    5469.17437290637, 5500, 5500, 5483.83673940805, 5360.36905140873, 
    5260.29028350104, 5143.41858983545, 5169.18439567109, 5257.74844319882, 
    5335.91671844887, 5395.07235242376, 5437.67757751002, 5474.19561320472, 
    5493.71445996705, 5430.26574678659, 5370.60392416211, 5299.05657156945, 
    5196.80336809989, 5069.26580954793, 4866.72364858187, 4550.00529703301, 
    4285.0086027095, 4006.44068169054, 3682.71566565236, 3791.61444283583, 
    4078.23388936473, 4351.05184542744, 4594.58757010561, 4722.15271796554, 
    4779.07571895829, 4807.87830856371, 4844.12526682691, 4880.78018042028, 
    4890.55569772915, 4871.10884857863, 4842.79479775391, 4784.69934096782, 
    4725.54558142431, 4650.47481124489, 4573.66469284064, 4520.29978028021, 
    4475.84585361604, 4426.7277390219, 4400.78026752467, 4388.60470794046, 
    4405.39850516058, 4419.18185522252, 4419.18185522252, 4391.36072790091, 
    4387.24020636153, 4361.18105035316, 4377.1518112124, 4399.48725672492, 
    4419.18185522252, 4434.06810454889, 4444.32257161226, 4462.33390411988, 
    4469.27439050223, 4478.96262991551, 4456.34441745014, 4408.25175552487, 
    4333.15956160189, 4276.47391966707, 4226.25248476706, 4193.88147434925, 
    4148.86631177499, 4102.41995330455, 4037.37862020813, 3967.01842774026, 
    3926.67892396058, 3911.01992262912, 3895.15734030234, 3868.82495086147, 
    3837.22582361098, 3807.9400935436, 3768.83194811735, 3708.48246321943, 
    3619.63273614653, 3499.54350243797, 3392.57529844592, 3295.30575471839, 
    3279.16880614892, 3301.29622115887, 3332.33277576082, 3328.19817106383, 
    3328.71685471083, 3287.97616131112, 3213.72721854304, 3114.97752235752, 
    3014.5461774317, 2898.91970776548, 2758.41088867188, 2592.33882768482, 
    2429.97449208961, 2080, 2213.26474854831, 2352.13760503619, 
    2664.28935020694, 2878.89007419664, 2941.06245126413, 2864.38591661102, 
    2659.74770600057, 2575.7707942982, 2576.24857471093, 2299.41904966201, 
    1627.01346544413, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 140, 888.509339995134, 
    1342.94244803009, 2075.11359247809, 2863.21289176457, 3499.27850908869, 
    3915.1221823787, 4073.9421829804, 4173.47329550756, 4207.47979745731, 
    4330.72884842842, 4405.36246428243, 4386.33120714808, 4294.20239844954, 
    4148.89562555905, 3951.59175146741, 3721.27612304688, 3485.19808803099, 
    3305.02901436926, 3239.79849281829, 3360.05065046364, 3569.89305986303, 
    3759.0490666634, 3935.98443056228, 4067.65515987029, 4164.81403268421, 
    4206.79498082343, 4195.10791681954, 4101.77248400289, 4108.0318649997, 
    4269.95679598799, 4538.45119423205, 4786.43706491839, 4920.06106739245, 
    4931.38438026846, 4864.50391133594, 4767.87269849225, 4632.48574314097, 
    4419.18185522252, 4134.69272413904, 3916.446095645, 3757.8187335117, 
    3662.63560900714, 3688.81729400881, 3790.7699812209, 3794.94622822043, 
    3768.14069260434, 3703.15717101759, 3611.44995937989, 3825.80800281077, 
    3943.22006109828, 3962.66125516521, 3881.13285731379, 3623.86417500358, 
    3237.10266690573, 2672.26131175894, 1986.93010261083, 1517.78682244505, 
    1280.12060546875, 1003.00093143071, 886.775249419965, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 2513.34521731361, 
    3088.95909212837, 3695.14468585039, 4307.41074153175, 4793.64067525731, 
    4968.77805804185, 5011.47023709696, 4955.62283052174, 4856.76331012619, 
    4711.72291358198, 4579.13970120788, 4420.81733847325, 4260.98641017652, 
    4008.0817335675, 3777.40123812498, 3540.37340362103, 3441.24200060235, 
    3425.80479829355, 3425.60405432324, 3496.41353104715, 3631.77664372094, 
    3826.6013490797, 3946.53839756857, 3804.35554060281, 3372.54430077798, 
    2603.84372784751, 2080.62891686437, 2398.75535520152, 2758.41088867188, 
    3241.21259093714, 3498.46508297279, 3736.5736263473, 3992.09927034817,
  4020.98003560274, 4110.87598049751, 4125.49551463753, 4145.25319183251, 
    4131.05399162064, 4096.30076991929, 4082.37446019618, 3973.29622277928, 
    3750.58816340872, 3493.90611879116, 3376.70554859439, 3495.91386246432, 
    3431.5629432299, 2793.98100974274, 2147.05598198693, 1526.58513556289, 
    -0, -0, 70, 70, 50, -0, -0, 50, 60, 70, 70, 70, 90, 150, 200, 
    274.994700677069, 370.154968261719, 370.154968261719, -0, -0, -0, -0, 
    1965.78910601674, 2709.90646152977, 3480.34565292378, 4046.04675631441, 
    4403.68854962397, 4360.7415958614, 3854.23560852992, 1766, 
    2806.41312168542, 3177.05319419266, 4127.60571680825, 4377.75052103451, 
    4377.75052103451, 4173.77830847508, 3934.42105296627, 3987.05075749315, 
    4300.63205301079, 4499.35434068869, 4537.85202096525, 4477.31624877846, 
    4326.74555073548, 4099.14472882657, 3753.54535048843, 3324.98107361783, 
    3314.11705486436, 3611.8971329163, 3950.97378862844, 4183.0489039971, 
    4222.17774212697, 4154.8172099826, 4147.18960648228, 4330.11179368499, 
    4362.73395111234, 4351.99607230612, 4154.29938028858, 3797.80523353718, 
    3469.85139461732, 3277.61142208088, 3212.34859573816, 3141.93719942548, 
    3263.62989777126, 3543.71394694577, 3733.72838607911, 3903.7209408581, 
    4163.15143546118, 4361.75548067696, 4489.32957678659, 4556.70929267321, 
    4549.09425735726, 4473.05960977483, 4318.99952864969, 4264.99278228124, 
    4194.82463765688, 4177.60458154242, 4148.40438854051, 4445.74677237223, 
    4805.08828117067, 5069.92798687305, 5333.47124508177, 5500, 5500, 5500, 
    5500, 5372.86910480702, 5242.74303103917, 5130.25233437584, 
    5166.54972835258, 5284.04435587133, 5383.9773433194, 5431.05300919888, 
    5475.86269708285, 5500, 5500, 5444.07720585174, 5358.0047742136, 
    5268.17305411743, 5143.41858983545, 4973.08800251612, 4707.14995191969, 
    4371.37063422808, 4076.50330509348, 3806.97997147211, 3608.34319408795, 
    3878.16869175898, 4125.21675734387, 4407.1378780158, 4645.54796870032, 
    4737.15944529165, 4812.41201955467, 4858.23537285806, 4902.12632099794, 
    4931.3626320052, 4921.11820393813, 4893.44118788322, 4888.422424769, 
    4861.98121897272, 4806.83587038517, 4729.98277396797, 4642.94767304985, 
    4577.32827821529, 4525.74384764616, 4478.09677073924, 4449.377366333, 
    4438.5461376554, 4445.19978724718, 4454.18758853827, 4450.07112799633, 
    4427.41478234726, 4399.69936778592, 4352.04903865383, 4369.08196953033, 
    4384.64155209726, 4399.46010685339, 4421.02593930867, 4424.65597379426, 
    4434.67276108499, 4439.12526963434, 4441.1709741073, 4419.18185522252, 
    4374.23018767839, 4306.16273464016, 4247.24746011692, 4210.92146191242, 
    4200.8162299973, 4167.19721586955, 4127.39118874191, 4068.26171991917, 
    3999.52398215101, 3954.46078736527, 3934.67776756083, 3915.74542323274, 
    3886.34229285979, 3851.64113706594, 3826.82067743905, 3788.32347940422, 
    3721.56627250762, 3629.56308221375, 3495.41460521863, 3387.2978515625, 
    3288.42038457, 3279.40182782013, 3314.38470408791, 3354.87379204938, 
    3358.54775809614, 3376.24288632733, 3353.62711448183, 3316.09664355681, 
    3245.44518255579, 3164.18490316693, 3072.46849956002, 2947.62370771738, 
    2780.95923433615, 2581.5445977205, 2350.38188836285, 2205.32990334674, 
    2237.18909749394, 2558.59012461617, 2803.93815541803, 2890.75420341085, 
    2871.38164711842, 1785, 2597.10589078815, 2647.60014105104, 
    2541.76195354153, 1824.39297967016, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 140, 315, 
    1280.9410291054, 1762.1339145278, 2429.75371674337, 3098.70357397284, 
    3632.32910174928, 3953.93321958808, 4043.53023923346, 4190.37634633393, 
    4266.25501340413, 4393.03079740587, 4449.32532201398, 4419.18185522252, 
    4307.91098703792, 4132.27451129727, 3923.02932270126, 3691.27712291416, 
    3451.31049769222, 3301.36392296107, 3304.95562032114, 3421.30003185411, 
    3639.45215542422, 3832.16463473204, 3990.32163035538, 4112.9578962823, 
    4194.32388560492, 4198.31337375572, 4145.80355055884, 3997.97899152185, 
    3924.14764711083, 4104.85956358721, 4446.45362578736, 4727.58474444727, 
    4904.33986470546, 4934.49487637794, 4879.56238600608, 4764.20403271419, 
    4576.17253522691, 4241.70944382539, 3943.01792879032, 3576.13967506267, 
    3264.90597502975, 3110.65078497658, 3166.75638153409, 3298.15943592975, 
    3358.83699334926, 3370.02645548351, 3208.71985883551, 2998.76333852398, 
    3168.52219272434, 3543.48806317734, 3692.87797799918, 3663.10655196715, 
    3387.2978515625, 2973.65730852926, 2279.85860533162, 1630.66287657026, 
    1281.01342162356, 1034.87945429264, 845.680345852758, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    2680.75179634465, 3474.51603522522, 4175.79852972415, 4723.49311933025, 
    4951.26098938805, 4982.57304229887, 4942.78876184155, 4831.24089860372, 
    4663.58676808772, 4511.51116016754, 4328.35890638688, 4142.15087633108, 
    3885.45323498966, 3663.38241160325, 3462.9457843413, 3472.99631161449, 
    3524.79863780112, 3575.00710815439, 3647.17702051727, 3748.66337242655, 
    3898.21047639002, 3980.55147725555, 3802.55183567699, 3334.71007829362, 
    2554.00631572143, 2051.66399533274, 2332.21304065897, 2628.07088373298, 
    3090.88041127282, 3318.99923275713, 3610.84804789616, 3866.32879320694,
  3874.08450079131, 3995.13176263748, 4045.10593260771, 4077.60900645708, 
    4086.16568765417, 4043.70136117229, 4033.38140758712, 3939.85575287349, 
    3734.25378737815, 3506.99108031804, 3405.36761594621, 3376.70554859439, 
    3274.43196168079, 2542.89508911879, 2032.992538224, 1383.69693130034, -0, 
    -0, 80, 80, 50, -0, -0, 50, 60, 70, 70, 80, 130, 210, 298.314826814311, 
    410.949909483355, 521.219387177922, 521.219387177922, -0, -0, -0, -0, -0, 
    2277.97651403559, 3082.76496174273, 3829.20900077229, 4194.54330180291, 
    4205.46200331951, 3850.37551549337, 2121, 3086.29108574574, 
    3643.31554328002, 4484.43366067841, 4689.25368557932, 4619.70235051738, 
    4343.14166107394, 4007.64152181727, 4065.89147763595, 4292.10229809536, 
    4498.83488353982, 4537.8222538012, 4460.48872867187, 4288.07212714434, 
    4065.89147763595, 3737.13173244481, 3372.33477803192, 3242.13974191054, 
    3497.56380949886, 3818.17171433262, 4040.96816153821, 4040.96816153821, 
    4012.3068596769, 3978.23737605758, 4163.30613282104, 4246.60980029448, 
    4259.93749761403, 4106.71828087391, 3765.09670526952, 3567.64221819272, 
    3405.54222609621, 3344.92609710997, 3279.49550040514, 3387.2978515625, 
    3657.27894794261, 3863.05374444867, 4036.22303570849, 4237.59973204695, 
    4432.00320790418, 4584.16237640955, 4630.53464153027, 4629.04910576852, 
    4516.04731594144, 4318.48556191764, 4251.44538670247, 4151.53502608605, 
    4176.57571639362, 4138.70106575482, 4531.64084091116, 4877.51731573073, 
    5133.05873194192, 5394.14176279953, 5500, 5500, 5500, 5500, 
    5369.02433461183, 5220.46377176872, 5130.25233437584, 5190.82614895916, 
    5329.83328664977, 5424.40173826285, 5475.83619567022, 5500, 5500, 5500, 
    5442.76209027326, 5328.09501231314, 5206.63588177411, 5041.90715228769, 
    4836.0688560959, 4524.08126839425, 4210.37300172984, 3835.87512321944, 
    3592.78905722457, 3656.04179032107, 3937.52422423681, 4189.92289850897, 
    4480.20313943056, 4671.69738551814, 4758.99827923559, 4840.22767163528, 
    4904.09066630066, 4954.66071893184, 4967.04911608482, 4944.23384052805, 
    4918.90422063861, 4917.11133839663, 4913.14148239435, 4886.93739508741, 
    4825.83335026585, 4737.09387160591, 4662.96766869414, 4597.31413723506, 
    4550.04507474109, 4520.2673219094, 4508.26971666312, 4500.72600227136, 
    4508.42513797794, 4489.99560003864, 4456.02663900666, 4419.18185522252, 
    4353.65551246436, 4355.93040511067, 4359.44735426831, 4377.57471234496, 
    4405.59926830213, 4402.4888231244, 4419.18185522252, 4423.44058553815, 
    4405.48493854552, 4363.20714934771, 4332.47754878125, 4276.05346605494, 
    4218.54580312429, 4193.01638850146, 4195.2688040095, 4182.42853355463, 
    4146.4752385024, 4091.1409456046, 4028.75710796791, 3980.26951185944, 
    3956.47104260958, 3932.7518404385, 3898.60027366041, 3861.05051401133, 
    3835.31157652327, 3799.17766028697, 3730.29412068192, 3634.03560632855, 
    3485.51506484745, 3367.50866370819, 3274.35469943958, 3277.03684312909, 
    3321.23393853857, 3387.2978515625, 3408.18782708944, 3433.42122945666, 
    3426.51116766018, 3404.6326325746, 3359.59776181611, 3300.91791950225, 
    3236.03268336836, 3138.37371030514, 2976.71698301131, 2758.41088867188, 
    2504.72405891937, 1785, 1650, 2445.83939218361, 2711.37703907259, 
    2826.30466735297, 2814.76949110804, 2743.70284981141, 2684.54737109843, 
    2692.27295204277, 2643.28529934411, 2015.67080270707, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 916.872621444644, 1296.29618994982, 1837.40155352749, 
    2264.38798679109, 2804.26705664742, 3327.40211292897, 3751.19910002766, 
    3996.05642896097, 4098.2137275811, 4300.97784669011, 4384.49354659516, 
    4468.97641542817, 4492.85745021801, 4444.94113327329, 4302.64777591844, 
    4115.61347479953, 3886.31023548027, 3668.84634131241, 3440.53381298654, 
    3310.69920417962, 3363.8337871381, 3505.40203139068, 3721.27612304688, 
    3908.93684160013, 4040.90067055146, 4150.98545849073, 4214.29882531785, 
    4179.66700157251, 4092.22175279345, 3894.53091252973, 3773.48969844624, 
    3907.30923731631, 4338.10272700369, 4677.4032198414, 4878.2126521227, 
    4926.96076597297, 4867.25824804016, 4712.32171919468, 4434.1763963412, 
    4065.89147763595, 3705.93311331032, 3257.56227907263, 2731.61080977136, 
    2698.18379410484, -0, 2875.96794095977, 2807.59814902013, 
    2831.39580724244, 2637.16488546979, 2578.04347065192, 2453.37220270061, 
    2922.53995945702, 3320.05933718933, 3348.03382908262, 3155.92683606048, 
    2696.4953142823, 1958.26070698089, 1441.60059236959, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 2373.87771358834, 3332.8622065098, 4065.89147763595, 
    4636.85794450593, 4936.12650235304, 4937.22251356404, 4929.07640290064, 
    4801.67484447686, 4610.68999242962, 4420.37730548988, 4195.13250407663, 
    3993.07296657111, 3736.87135620566, 3555.28486111031, 3449.00929133334, 
    3558.46627777804, 3668.42405108998, 3747.96983880879, 3810.2756154235, 
    3880.60496352852, 3975.63725055291, 4009.22748142413, 3793.2554891911, 
    3289.39729725054, 2532.0927203219, 2019.41089238274, 2283.72217145325, 
    2504.79604307267, 2914.34818667752, 3115.48068711273, 3455.57546519106, 
    3721.27612304688,
  3600.51660974093, 3754.36218200817, 3918.56507912478, 3981.07102017852, 
    4021.34943878696, 3999.43536104296, 3975.63113851771, 3894.95990373959, 
    3703.29958582433, 3473.60876600481, 3387.2978515625, 3349.88313888819, 
    3116.98776207318, 2349.67155892272, 1903.70624298749, -0, 0, 220, 220, 
    110, -0, -0, -0, 60, 60, 70, 70, 100, 170, 294.462890625, 
    454.557847665543, 630.451098056706, 762.080341837945, 845.523272431619, 
    845.523272431619, -0, -0, -0, -0, 1896.81606097386, 2524.51553257108, 
    3367.77049108889, 3836.14479047013, 3938.06268892357, 3710.7912185851, 
    2121, 3350.99352942098, 4285.86490557478, 4758.49111464245, 
    4984.58336246854, 4893.93022272587, 4525.63907762405, 4137.87163062236, 
    4148.87293797451, 4334.8991324368, 4476.17256113396, 4501.46585779971, 
    4391.61503501709, 4235.22510021712, 3981.73198172709, 3675.25671944374, 
    3372.33477803192, 3152.09306204873, 3358.45689206052, 3654.69630914649, 
    3808.7856062598, 3843.69126633846, 3771.81736295996, 3735.46645726738, 
    3885.97030478214, 4080.14136591005, 4154.3466437368, 4030.04168829123, 
    3633.74208681107, 3647.74954879378, 3555.50456295115, 3498.22448306192, 
    3460.63974664163, 3578.26645378281, 3825.08281353855, 4036.06030210206, 
    4219.43379573845, 4338.96597179017, 4535.45507253282, 4705.09398992894, 
    4741.48442926469, 4725.59197970421, 4522.47177777648, 4338.99003767761, 
    4153.68462542221, 4111.43922326499, 4150.47921499227, 4221.85947896899, 
    4606.81038385715, 4923.18099000978, 5198.27223244239, 5435.58585509719, 
    5500, 5500, 5500, 5500, 5349.85895251621, 5162.99428737976, 
    5125.71940048732, 5216.76360808599, 5385.52914519415, 5464.90301476158, 
    5500, 5500, 5500, 5500, 5405.74420495963, 5275.86410372662, 
    5121.68965739225, 4931.04948553095, 4687.47913753008, 4347.59768297222, 
    4004.43239823042, 3591.28159086951, 3500.09576918126, 3710.04738605745, 
    3985.38250808188, 4286.97957683877, 4546.80863170634, 4705.17867273803, 
    4792.70081294552, 4867.61249751165, 4938.96055982813, 4994.59804880115, 
    4993.68616805693, 4963.47509356863, 4932.75431889387, 4945.02112344743, 
    4964.33712908335, 4958.76507902168, 4915.39060701081, 4852.90512178117, 
    4781.80616572199, 4707.59059336081, 4665.47699760893, 4626.41681218195, 
    4607.89813696178, 4578.32663679459, 4567.08349472338, 4530.29954585172, 
    4483.18388534106, 4432.08885390189, 4369.84425878902, 4343.04028715643, 
    4346.5798099475, 4365.56415476479, 4397.05076590353, 4388.34263976385, 
    4399.09927684575, 4405.91823218844, 4373.01282338377, 4335.62153898393, 
    4290.77475823874, 4237.94784301508, 4179.68900127729, 4156.5010392446, 
    4157.04570439537, 4172.07565678349, 4149.93508416408, 4104.02761504217, 
    4043.54950615076, 4000.30916707978, 3976.17314769816, 3951.45314735884, 
    3908.2984315297, 3861.85068694359, 3832.11763325927, 3797.4173223791, 
    3730.47151565981, 3625.63420529593, 3468.50099902666, 3338.73312629021, 
    3252.13264817799, 3269.6989208843, 3328.01624230505, 3403.45813403919, 
    3452.29424454284, 3492.16198522141, 3507.07759271948, 3496.37125900719, 
    3466.50243893352, 3431.86034084497, 3396.49559766478, 3324.61713844296, 
    3181.94467214068, 2948.23263541471, 2663.12728238167, 2379.89224947935, 
    1785, 2345.62948429781, 2595.89799309203, 2693.9669471368, 
    2656.65718822161, 2643.48562327121, 2684.54737109843, 2701.74731743772, 
    2673.0796043214, 2154.2040825047, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 864.470906018281, 
    1282.13850005533, 1878.03207973945, 2437.220648202, 2824.62480659546, 
    3228.11091529902, 3587.50555599019, 3893.1433301861, 4065.89147763595, 
    4225.39353348885, 4406.49354238126, 4479.7056454309, 4528.79584731768, 
    4514.15358933247, 4451.63665279699, 4304.48459098614, 4122.97846447664, 
    3892.69040959579, 3684.77998399031, 3478.0847066637, 3387.2978515625, 
    3481.66253502784, 3641.16745293053, 3838.98566770243, 4009.50613461293, 
    4121.20790270203, 4211.39983449879, 4246.2876878849, 4198.00627762556, 
    4065.89147763595, 3827.83077691469, 3661.8414572119, 3755.99301464095, 
    4196.71842887763, 4625.14045090508, 4839.92667199204, 4898.93234642867, 
    4802.77141421831, 4537.1106517919, 4177.78207736749, 3827.04212989355, 
    3400.42013324701, 2823.83737196578, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    2302.97202081386, 2800.70871188519, 2934.94553825962, 2862.29063105759, 
    2364.65367009709, 1628.37549565869, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    3134.4535583085, 3973.57909249531, 4537.60774241509, 4909.95579886239, 
    4937.94684394875, 4903.8818839012, 4768.4691612025, 4569.52324865989, 
    4307.56064840759, 4044.10836611177, 3804.87336229593, 3583.72710852326, 
    3487.1683995268, 3515.76545611652, 3688.25682611362, 3849.32610431985, 
    3956.05809415576, 4008.1960916619, 4050.56696480522, 4081.45478883455, 
    4065.89147763595, 3797.50802943583, 3258.64385738585, 2492.43202030445, 
    2026.49670433428, 2247.067241975, 2393.17101842457, 2651.85719166634, 
    2817.45634588301, 3160.32060748104, 3431.09480450202,
  2962.79979085411, 3309.57716319209, 3793.86455577301, 3913.80502836861, 
    3955.21666608716, 3950.01759338794, 3921.55033721675, 3845.3996171513, 
    3679.30387576572, 3444.76981635978, 3312.74689984487, 3273.36570689209, 
    3005.87447990969, 2231.99400833569, 1796.81589981827, 1261.70589191854, 
    951.024886396472, 508.799507680931, 240.561416625977, 110, -0, -0, 0, 60, 
    60, 60, 70, 110, 210, 390.081193261582, 666.86758615337, 
    913.885148059206, 1030.12504413904, 1148.74554377555, 1148.74554377555, 
    878.370046558423, -0, -0, 100, 100, 2191.85384798669, 2711.0968746487, 
    3504.47209257673, 3628.66548190984, 3236.56938058759, -0, 
    3501.23942576116, 4751.26248240066, 4941.01607697947, 5084.13349441629, 
    5084.13349441629, 4722.59803316852, 4237.60231746056, 4148.47261273785, 
    4351.79388327314, 4427.33859517961, 4419.18185522252, 4301.47718662968, 
    4145.03316052522, 3923.77455605232, 3640.90782352977, 3350.74446580698, 
    3065.78548661781, 3248.36686089744, 3458.0544598461, 3535.98758921285, 
    3608.44980711514, 3527.86388672589, 3490.50886643424, 3547.54554998522, 
    3865.3906679157, 4026.49357584999, 3942.53929250717, 3691.62375259265, 
    3802.22636823206, 3756.77812986575, 3676.00657119448, 3561.66585465116, 
    3775.45161285051, 3998.65167303282, 4149.88950678816, 4374.06430209034, 
    4497.05297702495, 4660.88394442164, 4813.22280928466, 4850.28039058789, 
    4779.07571895829, 4524.60666365881, 4361.36170938685, 3873.16724161553, 
    4018.83518866473, 4018.83518866473, 4290.80718335442, 4600.38201967219, 
    4978.98548851565, 5230.73615401352, 5488.00621057352, 5500, 5500, 5500, 
    5500, 5297.94778862398, 5043.83854442317, 5100.14287797938, 
    5255.49434114642, 5453.4825529179, 5500, 5500, 5500, 5500, 5500, 
    5367.21422148121, 5218.58818763401, 5031.78736993824, 4841.08714239925, 
    4602.04179836577, 4276.34954295782, 3779.53635330664, 3442.32112419405, 
    3506.79123730342, 3791.56664398404, 4065.9990480495, 4371.87384428082, 
    4625.08393079456, 4764.92062851632, 4834.14237486198, 4892.49552853414, 
    4965.18281828652, 5020.62303800486, 5015.54520830443, 4970.61231682853, 
    4939.05947066118, 4959.04940587794, 5006.48837527728, 5012.58359123931, 
    4987.99494369202, 4937.99037066563, 4871.62972819122, 4814.29835567239, 
    4781.86020943425, 4739.21407877603, 4710.43115873538, 4654.93282205641, 
    4619.32391310962, 4563.85419120579, 4513.7246674622, 4460.7890428605, 
    4388.8528002745, 4360.6234774435, 4362.57585113177, 4379.31964194276, 
    4403.28829992248, 4401.06998914551, 4393.90218837798, 4388.61024663903, 
    4359.86130099612, 4329.04367736274, 4276.16524193238, 4214.60357565602, 
    4152.22008187518, 4120.04230865935, 4118.93192082208, 4148.7690733788, 
    4137.39600794016, 4104.5174815738, 4053.40615271908, 4013.4458781083, 
    3986.25537323231, 3955.04715247315, 3894.93874745134, 3844.00219279919, 
    3815.24315886467, 3791.71675268833, 3722.70509155187, 3608.02479336238, 
    3421.0003764866, 3311.23579024048, 3232.25130841111, 3260.75864248906, 
    3324.40770755227, 3409.74011133101, 3482.4642587378, 3521.06330496502, 
    3553.43380824945, 3555.12567695203, 3539.61844717339, 3510.27432203613, 
    3496.59114230658, 3449.59925950254, 3327.86111605462, 3133.93079348539, 
    2846.43522573809, 2538.83988991019, 2313.77075684498, 2050, 
    2417.69328328739, 2508.61798727007, 2546.7751121441, 2426.05821625029, 
    2684.0948877042, 2650.15288586886, 2673.7456790835, 2156.98066441291, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 0, 339.548167860464, 370.154968261719, 580.953491210938, 
    1045.44981682196, 1747.90439053496, 2501.39281145455, 2948.63036605486, 
    3291.77188105109, 3583.60737361876, 3798.60025079661, 4010.72000812187, 
    4157.30935116646, 4355.52383149408, 4480.58723664048, 4534.11677777774, 
    4541.55260432985, 4488.29899413952, 4435.39739488453, 4296.00473727452, 
    4129.37893206661, 3921.06932276618, 3708.74451889229, 3543.70356991625, 
    3507.21516882358, 3640.57524626332, 3804.95265992094, 3959.16279665329, 
    4102.24767120736, 4210.87364878938, 4257.27539539018, 4259.57711351582, 
    4208.33194106035, 4040.79093975107, 3798.56988909207, 3665.97085543583, 
    3728.12599853477, 4100.21024258561, 4582.4370534413, 4802.74048534601, 
    4850.85384233653, 4679.49038909916, 4321.02816131746, 3967.93812205799, 
    3551.30284304626, 3010.49242758443, 2269.3537644208, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 2309.32732346745, 2353.59573677407, 
    1959.99774656831, 1314.03726861552, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    2788.53514152859, 3853.42804331067, 4467.53877501883, 4877.45163932016, 
    4962.60360150187, 4847.82007699477, 4726.78813205612, 4484.98888794377, 
    4217.85417865135, 3921.93432647282, 3648.39858581575, 3468.59378580683, 
    3468.36100990915, 3623.80264473391, 3843.86633582009, 4029.02287517157, 
    4137.07116796901, 4189.07980354225, 4204.78239547505, 4198.7632260923, 
    4142.04472220311, 3807.46426300412, 3255.42143705721, 2448.4551413522, 
    2038.35750830864, 2246.71871222056, 2273.17799143101, 2423.09123895168, 
    2567.24792310544, 2828.38414264501, 3010.48588380405,
  -0, -0, 3693.47392053245, 3843.41483075604, 3893.0976069997, 
    3888.5919653795, 3858.06099281311, 3797.72737991075, 3672.28208036543, 
    3410.1662854819, 3170.69713917441, 3202.46258709802, 3045.81887857155, 
    1990.6807815108, 1773.40783977158, 1320.4348340318, 1022.21679378907, 
    594.35588556263, 240.561416625977, 110, -0, -0, 50, 60, 60, 60, 60, 110, 
    240.561416625977, 568.129851826152, 988.534416165442, 1269.72442032015, 
    1295.45252832193, 1539.40042009849, 1642.90993477833, 914.096642193625, 
    -0, -0, 100, 100, 100, 2075.60747320127, 2932.05165249865, 
    2932.05165249865, -0, -0, 3430.46696330043, 5329.45434438846, 
    5205.16097458755, 5427.23443154278, 5256.74918021299, 4905.86657626604, 
    4375.36302753054, 4008.88235563241, 4351.79388327314, 4352.73119834405, 
    4305.28875358758, 4178.17510452637, 3979.21947176779, 3830.11702609303, 
    3578.60201942324, 3277.04056783429, 2852.34067351616, 3013.92259237114, 
    3259.79219657543, 3324.96684274053, 3324.96684274053, 3302.92837298805, 
    3263.36088012671, 3202.78218182126, 3796.50696862539, 3933.81447138312, 
    3841.30589825508, 3863.50694751772, 4017.67660052303, 4017.67660052303, 
    3993.66484555998, 3755.77009628042, 3907.96679995516, 4187.07201531878, 
    4317.1441062516, 4540.31970083137, 4655.97848076932, 4793.57375813843, 
    4910.50591563576, 4935.31973389305, 4791.54877792303, 4596.3672340807, 
    4393.99069254706, 3919.58454510099, 4018.83518866473, 4023.35797557429, 
    4307.90604945332, 4721.04219163916, 5080.00878239453, 5149.62846344049, 
    5500, 5500, 5500, 5500, 5500, 5337.74846622265, 4804.99364610812, 
    4940.24179224618, 5318.07171213997, 5500, 5500, 5500, 5500, 5500, 
    5488.90083218743, 5321.29224917016, 5125.89485568776, 4938.14519554415, 
    4836.37486225826, 4603.19767756157, 4300.29602119776, 3447.09075757024, 
    3275.44737597374, 3587.38967313604, 3886.11670221938, 4092.03298882453, 
    4388.72723864802, 4718.27732420735, 4856.8715877509, 4873.21101694887, 
    4932.47095827107, 5016.23281999194, 5076.45471014727, 5052.08322456832, 
    4933.65535947585, 4898.51392502816, 4948.71364982782, 5050.66235575904, 
    5055.73466537868, 5055.14029294882, 5018.35572117712, 4963.59185600792, 
    4933.21533256016, 4902.34340319053, 4847.45281878129, 4809.37357072554, 
    4728.43034004637, 4670.89129103325, 4621.14999850827, 4546.4587792182, 
    4513.33703257819, 4441.97893410865, 4419.18185522252, 4433.13845946233, 
    4419.18185522252, 4428.63953640388, 4428.04752570937, 4404.20797677294, 
    4361.16458442804, 4361.4594567772, 4355.04006535089, 4279.85243490505, 
    4212.09022014818, 4123.73282383519, 4065.89147763595, 4072.23904987904, 
    4117.21611961442, 4113.56145161891, 4102.61093948743, 4048.79356457996, 
    4015.48843245652, 3987.54320775852, 3963.58006214986, 3810.50780070054, 
    3783.38702789383, 3788.96450964009, 3779.15884088653, 3705.7667113168, 
    3591.26694701963, 3415.97309259398, 3289.49604039946, 3188.16819560817, 
    3258.79463837935, 3333.47906123188, 3417.99906966229, 3500.27971762395, 
    3549.89079093654, 3601.05561841165, 3605.48557779816, 3591.59957755486, 
    3564.5977815243, 3548.14993149421, 3553.78904390946, 3468.85940008278, 
    3317.4742980548, 3065.78548661781, 2795.95298181886, 2471.42213665709, 
    2216.39398385516, 1785, 2298.09772648498, 2412.09042801985, 
    2132.01586273906, 2595.75081203887, 2664.46510021082, 2650.15288586886, 
    1554.90424178863, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 0, 471.187348308304, 460.55078275968, 
    523.590127535382, 762.513365295387, 1280.30260554673, 2505.58449328403, 
    3122.39383096092, 3496.821383127, 3734.78057049221, 3915.40737035201, 
    4038.15973505623, 4186.29194690078, 4355.58440297382, 4490.87576645187, 
    4526.5136905016, 4573.65983921642, 4529.20334114466, 4459.19423354154, 
    4425.17146704128, 4269.77412505828, 4139.24202503657, 3946.17818963246, 
    3732.87245339223, 3622.42902701333, 3710.21265635764, 3831.20153441616, 
    3985.11168002264, 4087.33282808591, 4246.69801075964, 4347.00011927591, 
    4376.37378087523, 4312.10972391684, 4234.12437195996, 4035.39265904635, 
    3694.63556472288, 3670.39419970152, 3722.04431683386, 4042.11299462112, 
    4549.06325010232, 4736.928366173, 4737.84563344613, 4451.63842905357, 
    4111.12903024681, 3683.59740448296, 3137.06445755147, 2134.86566706509, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 2133.86241585732, 3484.58980582209, 
    4475.8117904227, 4844.68949305607, 4973.84937734333, 4762.04048977422, 
    4723.17706527218, 4384.29060121212, 4098.70152758828, 3796.5051380574, 
    3456.12211237543, 3387.2978515625, 3516.94966762434, 3747.78774189978, 
    4037.32803042488, 4218.26140353344, 4345.79663943338, 4360.24806104594, 
    4369.40275863863, 4307.18810144844, 4274.08924023662, 3872.95047162102, 
    3387.2978515625, 2295.82884100718, 2045.69272393484, 2150.79456281612, 
    2150.79456281612, 2149.90603733489, 2248.1157574043, 2314.74288836357, 
    2314.74288836357,
  -0, -0, 3554.34777004244, 3769.78737242693, 3832.13891521313, 
    3831.71425991423, 3805.99025284234, 3744.87559562634, 3619.40391795924, 
    3429.63864009214, 3184.48813854546, 3125.86567781183, 2841.08863476065, 
    1818.56640632364, 1881.14060203725, 1390.05342789468, 1004.75177194821, 
    602.981580668048, 240.561416625977, 110, -0, 50, 50, 60, 60, 50, 60, 120, 
    294.462890625, 726.308092174743, 1197.06655750824, 1463.47249798371, 
    1569.11829824086, 1564.83308930488, 1564.83308930488, 1280.12060546875, 
    761.027380776171, 100, 100, 100, 100, 100, 2164.02773492811, 
    2164.02773492811, -0, -0, 3271.71775086074, 5440.20634452369, 
    5339.64400063554, 5485.3823968402, 5354.91480193788, 4903.93892301634, 
    4493.21886751058, 4046.52921787512, 4008.85145397218, 4117.45108713962, 
    4301.69685564358, 4100.48465221441, 3796.55214795494, 3538.98062618728, 
    3368.27467074881, 3095.41683266998, 3102.37441254567, 3040.3200331431, 
    3040.10956882593, 3040.10956882593, 2935.11540877342, 2950.24941306784, 
    2968.70443710968, 3096.63266147184, 3555.95934908073, 3555.95934908073, 
    3579.46693947197, 4106.08911354369, 4224.11319180792, 4138.42121005116, 
    4248.35850551692, 4019.64671961504, 3958.29906111687, 4419.18185522252, 
    4526.97702858981, 4602.17388789255, 4673.35347529601, 4866.85089001879, 
    4948.15517064942, 4938.08053185085, 4760.53772990439, 4544.97853613992, 
    4146.70027563375, 4032.72565237008, 4024.36262100738, 3650.83489295673, 
    4319.63800020722, 4823.00011110016, 5123.70771464257, 5248.14481661078, 
    5500, 5500, 5500, 5500, 5500, 5404.39709258613, 4821.58211231518, 
    4782.95432082715, 5347.32619235432, 5500, 5500, 5500, 5500, 5500, 
    5441.21030767324, 5247.09444137839, 5034.39299332481, 4954.37624018006, 
    4826.81999416826, 4605.66375294979, 4298.96554699309, 3832.19776974225, 
    3503.32199654759, 3703.24884652643, 4041.43827120829, 4323.79252307969, 
    4572.12324659915, 4816.74087910556, 4941.78186814098, 4928.65839609328, 
    5015.61742186706, 5093.52340912613, 5098.69284361201, 5041.10994338398, 
    4913.2614841817, 4900.20402280406, 4985.91106986883, 5075.22056863895, 
    5083.84645364331, 5078.43366534473, 5050.80969206908, 5046.71667120691, 
    5004.02251548812, 4982.84544449888, 4933.69275593722, 4857.00905805189, 
    4766.41036453591, 4697.97564964142, 4662.45728409252, 4629.65878271456, 
    4581.56339876016, 4577.28389125153, 4549.57390311302, 4556.36932713984, 
    4495.57053185794, 4496.44341019521, 4467.4601066783, 4427.54326966898, 
    4423.24209503253, 4379.00985259985, 4371.16240301698, 4281.05344632322, 
    4226.43355911789, 4134.9264695589, 4065.89147763595, 4076.88850009272, 
    4066.81951874132, 4071.46197160478, 4065.89147763595, 4040.11887620579, 
    3987.13594637445, 3951.35930209838, 3933.10642495035, 3844.21620724753, 
    3782.60204554479, 3763.30905705176, 3745.63823852308, 3668.34315493024, 
    3546.711495913, 3387.2978515625, 3255.50354974473, 3174.26713700778, 
    3255.51795417638, 3349.4397680322, 3436.55484547946, 3521.60192231363, 
    3560.28465421395, 3605.42823366385, 3634.61522020593, 3618.29428726984, 
    3598.1374065553, 3563.89618587507, 3570.8093226744, 3505.33038509642, 
    3392.13403804304, 3213.78256696395, 2968.56659308582, 2676.92419493517, 
    2302.76783036108, 1655, 1979.21790283071, 1979.21790283071, 
    1739.35099441285, 2026.58477017108, 2269.52905210909, 2269.52905210909, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 60, 613.659905704199, 759.628478342875, 823.987360332972, 
    884.78125186968, 1137.36424270363, 1847.34841270392, 3048.32941115572, 
    3550.68408962737, 3877.26426803577, 4053.4957192982, 4139.60843570652, 
    4227.74279399881, 4336.11651902156, 4465.41350879073, 4578.85464533158, 
    4543.89573538835, 4533.41653866305, 4448.61669519406, 4339.94936898845, 
    4248.46311882686, 4208.34591689366, 4090.78699051155, 4014.59173670115, 
    3892.52694658128, 3877.45305313963, 3993.12361888003, 4102.45777477942, 
    4166.17727536142, 4275.70826398458, 4389.1560133734, 4429.44973777614, 
    4474.41101001641, 4444.78613091794, 4354.8200507453, 4065.89147763595, 
    3815.48894896475, 3598.01292515549, 3834.04476341042, 4118.19800200101, 
    4466.64350438487, 4567.34034510157, 4447.40460758244, 4081.46959759635, 
    3654.68434141869, 2952.65322169732, 2224.64586479383, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 1852.63707462624, 3307.2746589306, 4383.35526440598, 
    4731.30038550363, 4928.08078628642, 4863.21928864987, 4619.97150575679, 
    4344.68547530654, 3977.88389331053, 3691.09049396435, 3442.32155868052, 
    3398.81783013477, 3594.64417365018, 3899.94843274914, 4150.98574664692, 
    4341.96927252705, 4459.06281578567, 4452.86646435831, 4469.49580900383, 
    4448.97164021662, 4329.82978243286, 3923.06500019969, 3399.78889100431, 
    2376.61964955045, 2177.26284341851, 2158.13030892266, 2031.55280436304, 
    1898.57764014, 1699.69467065787, 1849.13407606054, 1849.13407606054,
  -0, -0, 3397.44401810969, 3698.66708000154, 3766.91236330139, 
    3775.55387986501, 3743.16985503757, 3673.56013080887, 3555.48168463885, 
    3417.04933227768, 3168.27094324108, 2950.05667639655, 2440.73259955919, 
    1897.08962201497, 1853.13515713095, 1447.31926549413, 997.022691148318, 
    623.086892222538, 240.561416625977, -0, 0, 60, 60, 50, 50, 50, 50, 150, 
    370.154968261719, 757.62064017006, 1217.64363692565, 1521.64019121917, 
    1668.34213770749, 1668.34213770749, 1626.85622178864, 1564.66624447886, 
    1102.91886923426, 100, 100, 100, 100, 100, -0, -0, -0, -0, -0, 
    5306.24355070167, 5425.30103647078, 5500, 5398.43095160084, 
    5038.42931731113, 4647.1419524814, 4315.86276734277, 3874.65748222161, 
    3953.66734382422, 3953.66734382422, 3976.66375494097, 3630.54826892853, 
    3353.09250015558, 3190.04968060018, 3074.31665359863, 3073.66777772667, 
    2990.75785186406, 3034.51703954189, 2959.36533400998, 2793.39347261145, 
    2650.07769064198, 2731.26883150826, 3041.28954690429, 3575.06898452834, 
    3657.30384960308, 4002.75377736383, 4276.97934675011, 4302.39016468742, 
    4292.33220250706, 4486.71510691601, 4458.06255843815, 4488.7296769409, 
    4546.28430499833, 4526.3804493744, 4537.40491236491, 4674.09104709944, 
    4828.64744133388, 4915.83428691809, 4848.02281725176, 4654.50349915327, 
    4341.71768164163, 3872.90000765855, 3851.1550854153, 3898.23542898295, 
    4040.04269753474, 4507.44464934351, 4857.98424897526, 5143.41858983545, 
    5194.96002699302, 5384.17823902997, 5500, 5500, 5500, 5500, 
    5483.45092270085, 5180.56518851386, 5062.26059618368, 5395.23886237639, 
    5500, 5500, 5500, 5500, 5414.59540251387, 5301.47302105666, 
    5174.03056390936, 5063.61714975878, 4919.86542151935, 4736.75309416276, 
    4527.52966199042, 4241.58826868122, 4068.19683615106, 3910.65757645228, 
    4000.1678814618, 4205.39764283441, 4446.70692819957, 4668.32830856867, 
    4888.82024772198, 5009.59918050319, 5038.07991041379, 5068.75685151982, 
    5082.00050165247, 5067.6408263323, 5024.23155752401, 4954.45106378305, 
    4973.95572771757, 5041.68454997079, 5098.4078684007, 5114.17818709175, 
    5108.81350745713, 5091.65029030573, 5077.86433086452, 5059.87022250982, 
    5024.96006291183, 4971.63891369344, 4896.19516857626, 4804.65267603405, 
    4738.38629163435, 4704.95524534954, 4694.02650063298, 4689.29677570612, 
    4693.42488442922, 4685.28520301608, 4648.66857823006, 4580.97403141904, 
    4545.37389309014, 4504.23592387839, 4473.02842275389, 4455.38663381978, 
    4420.40881182117, 4388.0400749683, 4336.50055889717, 4256.7069403626, 
    4161.40757914727, 4100.73612111718, 4077.6233310068, 4054.56433925547, 
    4054.56433925547, 4022.47183116564, 4001.77517858455, 3935.60410695724, 
    3916.25311383863, 3863.17879642857, 3809.33392509591, 3764.78069406236, 
    3721.27612304688, 3667.27566817528, 3579.21912315862, 3456.0633073862, 
    3320.64747912574, 3219.49179593401, 3195.02970490662, 3275.90429629344, 
    3371.18090417339, 3482.5835499255, 3573.14868531632, 3619.56649255178, 
    3643.56396371496, 3653.54325149758, 3634.41312376682, 3616.20522296175, 
    3587.76639908558, 3562.93010176749, 3502.22858114923, 3415.21695463938, 
    3282.12432243219, 3049.70892999427, 2740.07437723829, 2360.610379805, 
    1987.40516627892, 1420, 1420, 1420, -0, 170, 170, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 781.876492323839, 
    1101.54602050781, 1377.47256082051, 1519.47516769191, 1531.03090604792, 
    1838.65772747425, 2529.24000522928, 3387.2978515625, 3894.46463281704, 
    4191.26402076102, 4288.81831285344, 4337.33692850565, 4402.10011164659, 
    4471.86716201908, 4533.57235300289, 4561.13704570939, 4536.67913862573, 
    4419.18185522252, 4287.4288954186, 4201.73771297807, 4129.15178276053, 
    4112.73805502854, 4135.31413048706, 4148.56380480288, 4161.61132441949, 
    4233.19039674449, 4306.23584405356, 4399.3772951002, 4462.58780736448, 
    4545.25639319114, 4619.32438128673, 4658.26889089545, 4683.69418917165, 
    4647.96516619846, 4543.0351045128, 4340.91555500501, 4099.90082940081, 
    3839.39995688406, 3925.4371155894, 4136.98307315159, 4265.58753185458, 
    4228.81490905139, 3931.09536164217, 3516.05637332887, 2914.0450728526, 
    2128.80506391338, 1865.52205308119, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    3148.34353683309, 4132.700631571, 4544.19380268536, 4803.6962562786, 
    4779.07571895829, 4472.50680299603, 4222.70383627429, 3883.2278232621, 
    3589.69890500286, 3461.02104294905, 3565.64799467961, 3767.18515201678, 
    4040.60285518513, 4272.86768639955, 4419.18185522252, 4504.0114045564, 
    4527.71510091716, 4527.35126326417, 4482.04556947909, 4327.42370451067, 
    3905.82340479115, 3311.03200322251, 2588.87892345992, 2269.36128520721, 
    2158.13030892266, 1935.05359591651, 1651.95675953546, 1330.71650579107, 
    1537.3115201537, 1559.16208581883,
  -0, 2388.57623675491, 3367.85281415744, 3619.66239663698, 3709.87864513923, 
    3709.87864513923, 3674.58952291853, 3612.75529651687, 3516.50011147575, 
    3375.79613880516, 3129.26458720502, 2865.32456136072, 2191.85384798669, 
    1913.92108310739, 1913.92108310739, 1595.68136094379, 1027.05633797533, 
    581.449841399923, -0, -0, 60, 60, 60, 50, 40, 40, 50, 150, 
    402.475921288518, 857.046932314587, 1342.15366033827, 1682.53479734835, 
    1668.34213770749, 1863.68921468779, 1728.77993307367, 1605.25764654014, 
    1299.54956546752, -0, 100, 100, 100, 100, 100, -0, -0, -0, 
    2612.67595193276, 5326.5695224148, 5500, 5500, 5500, 5270.16008827164, 
    4816.77699305425, 4486.56528882751, 3965.96890536864, 3975.16045940429, 
    3861.25724741713, 3730.81399980191, 3617.02344207622, 3360.51271550433, 
    3262.57316863858, 3182.18907151254, 3099.42381208569, 3163.14284599432, 
    3180.42631254478, 3013.79914357568, 3001.96553694285, 2850.5906142414, 
    2735.5567231953, 3238.29484895795, 3639.77990372877, 3865.51998766253, 
    4009.23872192719, 4588.84627364909, 4656.87693236954, 4736.99993172626, 
    4757.88643930665, 4756.36445998903, 4760.64468068626, 4700.56084219836, 
    4508.53024717935, 4483.16938858982, 4565.68471984985, 4760.19446805797, 
    4760.19446805797, 4726.16010850083, 4472.73163722239, 4088.11748700698, 
    3944.30504466729, 3875.92853271663, 3851.74758236934, 4099.62581069767, 
    4611.15811463755, 4940.52495850275, 5195.74235543429, 5261.27543602944, 
    5365.38484636588, 5500, 5500, 5500, 5500, 5500, 5420.97277336356, 
    5322.58034781705, 5500, 5500, 5500, 5500, 5417.00006216016, 
    5266.229737004, 5133.4082546616, 5068.39528599829, 5003.38084314214, 
    4847.90850018906, 4689.11845084485, 4452.78559779699, 4319.86870400142, 
    4215.16094125673, 4248.06253426163, 4268.25993063181, 4347.78743847826, 
    4576.19651944405, 4785.52417478852, 4986.40730269058, 5089.36831849449, 
    5100.42616667328, 5101.98034069695, 5100.82618755528, 5086.70362149859, 
    5028.31731041222, 4991.92007143827, 5036.97973878683, 5099.51026057288, 
    5143.41858983545, 5150.9018023161, 5129.82225444412, 5116.1668351328, 
    5098.7687928, 5083.59398231801, 5044.99244153363, 4992.0657024142, 
    4918.38568205532, 4837.11864555884, 4779.07571895829, 4751.20318225928, 
    4762.80753793827, 4782.02731554737, 4787.57546359392, 4790.95225554494, 
    4750.62291039043, 4668.85848216747, 4606.78554948697, 4555.5735677832, 
    4520.68911497314, 4502.92379314328, 4477.15490319852, 4431.27367810259, 
    4374.5376444139, 4291.06117206126, 4209.32073079428, 4132.3485376696, 
    4084.7938622235, 4047.48960494793, 4030.06534627049, 3995.64058866003, 
    3974.81562459994, 3910.48631769647, 3881.15475247488, 3801.47181496258, 
    3771.48418179553, 3708.15329097954, 3637.41814960349, 3585.9080472431, 
    3484.21400137198, 3362.27162120994, 3231.83974259164, 3179.28728534177, 
    3213.4278166885, 3309.98728352354, 3412.06122897324, 3549.45359006281, 
    3656.30414949698, 3698.51190713644, 3707.18693868728, 3687.07734133377, 
    3654.88689803144, 3624.59401759438, 3604.97159702923, 3578.80803228658, 
    3512.74965776996, 3445.14305486669, 3341.98671451703, 3101.78992410471, 
    2787.86197977078, 2421.49228890813, 1942.97725485398, 1420, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 0, 110, 1138.005006741, 1632.53004636499, 2005.75717856688, 
    2163.51277666546, 2169.11125537514, 2510.41927870122, 3288.5626610895, 
    3930.46450430189, 4292.07083685926, 4453.71526367773, 4492.66735563317, 
    4518.44225208882, 4552.23600325462, 4582.76531271492, 4604.22503389036, 
    4549.30204363284, 4435.68730247372, 4251.53185423542, 4067.63492290258, 
    3987.54009933735, 4036.31068853482, 4137.66551680815, 4224.95495767824, 
    4336.73467898964, 4421.19929710537, 4526.74571961149, 4598.77075037642, 
    4670.66182545693, 4734.29342023652, 4787.44564447521, 4842.4847522657, 
    4880.8529608905, 4872.31795113008, 4839.94977248983, 4747.17541307318, 
    4562.2900566437, 4356.26226788742, 4110.07744630676, 4050.28750283642, 
    4128.06592859016, 4076.85031706946, 3794.26814264363, 3321.62006333797, 
    2885.79958513901, 2156.35015946004, 1527.80671560025, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 2772.18713919472, 3804.28055866373, 4372.42579560667, 
    4605.61216236217, 4654.91131060669, 4360.81854700825, 4102.2778035788, 
    3792.36201350218, 3538.30617355357, 3528.28000583467, 3706.23909232665, 
    3960.0784049736, 4188.56367548649, 4375.89911551203, 4467.49539121234, 
    4517.56979738172, 4552.36830289084, 4553.22102228948, 4515.20282617647, 
    4356.36025352067, 3913.10305022652, 3285.97138183125, 2604.25348161994, 
    2255.60286943255, 2121.33481741772, 1748.73555450518, 1340.30780384297, 
    -0, 1050, 1050,
  -0, 2554.6, 3332.7, 3586.3, 3663.4, 3644.1, 3605.8, 3549.7, 3469.7, 3339.1, 
    3065.78540039062, 2710.3, 2006.9, 1982, 1948.1, 1680.2, 1101.54602050781, 
    581.2, -0, -0, 60, 60, 60, 50, 40, 0, 50, 110, 433.2, 986.2, 1582.7, 
    1948.8, 1997.4, 2096.8, 1908.3, 1687, 1400.7, 0, 100, 100, 100, 100, 100, 
    100, 0, -0, 3452.9, 5500, 5500, 5500, 5500, 5500, 5082.7, 4681.6, 4164.6, 
    4078.7, 4037.8, 3873, 3809.3, 3451.8, 3324.9, 3371.4, 3486.2, 3609.4, 
    3618, 3445.4, 3441.8, 3363, 3373.8, 3818.5, 4158.1, 4384, 4511.2, 4903.1, 
    4953.8, 4987.5, 4971.7, 4958.2, 4906.1, 4792.8, 4455.3, 4386.8, 
    4419.181640625, 4631.1, 4654.6, 4504.2, 4198.9, 3947.8, 3896.1, 3767.9, 
    3892.2, 4249.3, 4717.8, 5049.3, 5261.4, 5310.1, 5378.3, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5273.4, 5132.2, 5004.8, 
    5007.1, 4932, 4784.1, 4572.4, 4423.9, 4375.7, 4379.9, 4448.1, 4489.3, 
    4509.9, 4677.6, 4885.6, 5050.8, 5127.9, 5129.6, 5122.7, 5122.1, 5103.3, 
    5061, 5059.2, 5097.2, 5145.2, 5167.7, 5164.3, 5143.41845703125, 5121.2, 
    5095.6, 5073.4, 5029.1, 4977.8, 4915.5, 4853.1, 4815.3, 4798.6, 4809.5, 
    4827.7, 4840.1, 4838.8, 4790.3, 4713.4, 4649.3, 4604.3, 4570.4, 4547.5, 
    4514, 4468, 4419.181640625, 4330, 4249.9, 4184.4, 4136.9, 4090.9, 4048, 
    4003.5, 3960.3, 3886.6, 3843.4, 3746.4, 3701.3, 3637.7, 3566.6, 3525.1, 
    3436.2, 3318.9, 3195.5, 3176.7, 3236, 3348.6, 3466.1, 3604.2, 3721.4, 
    3776.5, 3779.2, 3751.3, 3721.27612304688, 3676.4, 3646.1, 3613.4, 3557.6, 
    3473.3, 3293, 3065.78540039062, 2775.7, 2271.4, 1489.94085357879, -0, -0, 
    -0, -0, -0, -0, 253.361404418945, 253.361404418945, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 60, 617.9, 1537, 2120.4, 2554.2, 
    2795.9, 2902.2, 3253.8, 3812, 4272.3, 4521.7, 4609.6, 4616.9, 4624.2, 
    4619.7, 4602.1, 4556.2, 4445.3, 4306.8, 4128.4, 3987.3, 3996.3, 4101.5, 
    4241.3, 4391.9, 4546.2, 4660.8, 4779.07568359375, 4838.2, 4895.7, 4947.6, 
    4990.3, 5024.5, 5038.7, 5019.8, 4980.5, 4904.3, 4747.4, 4547.1, 4326.6, 
    4222.4, 4124.1, 3787.3, 3169.7, 2556.9, 2055.9, 1269.8, 150, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 3216.5, 3993.2, 4276.8, 4276.8, 4213.4, 
    3994.3, 3740, 3615.8, 3693.2, 3871.8, 4104.9, 4278, 4397.5, 4457.3, 
    4489.1, 4515.1, 4523, 4489.4, 4303.6, 3850.9, 3185.2, 2507, 2139.4, 
    2028.2, 1522.7, 120, -0, 150, 150,
  1569.41248786985, 2720.58896521007, 3297.6275131904, 3552.90195559347, 
    3616.86457611774, 3578.22265089216, 3536.93180511499, 3486.64163735172, 
    3422.90412364993, 3302.35500499044, 2986.55850596432, 2555.19959604575, 
    1822.02749545516, 2050.11157763661, 1982.33615119378, 1764.80571352535, 
    1156.20384022787, 580.953491210938, -0, 60, 60, 60, 60, 40, 40, -0, 40, 
    70, 463.933091178488, 1086.87921984415, 1823.20262702432, 
    2215.01638749791, 2326.42088691749, 2329.84780583561, 2087.89843681754, 
    1768.74629726939, 1501.84006182986, 1260.26187003645, -0, 100, 100, 100, 
    100, 100, 0, 2387.05420861712, 4293.19861384892, 5434.98257365275, 5500, 
    5500, 5500, 5500, 5348.69203814715, 4876.70711901058, 4363.1857579731, 
    4182.25942845203, 4214.41266049382, 4015.12379332166, 4001.65156057947, 
    3543.0419718513, 3387.2978515625, 3560.59406913485, 3872.97333251224, 
    4055.59693064124, 4055.59693064124, 3877.01434748693, 3881.69140743309, 
    3875.41865099034, 4012.0517591003, 4398.67290510145, 4676.51546230655, 
    4902.57319501789, 5013.23653260795, 5217.44823133, 5250.7021775735, 
    5238.04520011307, 5185.43374390872, 5159.99411426561, 5051.50012032997, 
    4884.97018924588, 4402.06387071145, 4290.38733174658, 4272.09849701926, 
    4501.91435261144, 4549.00365634982, 4282.14290184192, 3925.13659581978, 
    3807.41238367895, 3847.967479711, 3659.87962070414, 3932.68760983837, 
    4398.94795873548, 4824.41831283757, 5158.09963789504, 5327.14369041358, 
    5358.82825201454, 5391.14228077592, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5479.21252054366, 5129.77760708091, 
    4998.1719880531, 4876.10926941463, 4945.82061307843, 4860.71245222423, 
    4720.29403299393, 4455.65345146027, 4395.03800471817, 4431.59443408217, 
    4544.5545352906, 4648.10773574965, 4710.36866488924, 4671.96258966656, 
    4779.08832509019, 4985.72050885708, 5115.25005753508, 5166.51369512106, 
    5158.68120874739, 5143.41858983545, 5143.41858983545, 5119.84793338933, 
    5093.74714665131, 5126.42310942176, 5157.51065223425, 5190.94447492074, 
    5192.01768033413, 5177.72068086629, 5153.06559766094, 5126.13320011889, 
    5092.34639220261, 5063.11332266054, 5013.13781546362, 4963.50725387061, 
    4912.63341219333, 4869.01207643555, 4851.59958342481, 4845.97791298006, 
    4856.18203363976, 4873.37292940396, 4892.6073660056, 4886.73960387143, 
    4830.00320293584, 4757.98618227015, 4691.82218010777, 4652.97135655292, 
    4620.20300974627, 4592.03114347584, 4550.90860421466, 4504.7134311844, 
    4444.11049912336, 4369.02119211921, 4290.39442626971, 4236.38290837277, 
    4189.02521931735, 4134.40495570156, 4065.89147763595, 4011.42729298962, 
    3945.70668407593, 3862.67953999014, 3805.72952449419, 3691.40330968253, 
    3631.02577008132, 3567.27914023669, 3495.880473166, 3464.26871465791, 
    3388.13448812137, 3275.49543321328, 3159.14725230155, 3174.07742446859, 
    3258.61327059503, 3376.17978770714, 3520.21770714033, 3658.88860573886, 
    3786.55014589823, 3854.58070858104, 3851.30257095843, 3815.44291499685, 
    3776.26007491692, 3728.194576495, 3687.2261306164, 3648.09155770698, 
    3602.49041530468, 3501.50662670867, 3244.08098569645, 3026.60394967445, 
    2763.59213210414, 2121.22132124245, -0, -0, 1450.39623001455, 
    1806.10087615306, 1889.71053412127, -0, 1910.10809647039, 
    1910.10809647039, 1810.28645405115, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 637.728619557105, 1125.81390596563, 
    1935.96005823437, 2608.27121658887, 3102.56829594886, 3428.33327862068, 
    3635.27219323796, 3997.14469990194, 4335.44293546522, 4614.09777081994, 
    4751.24423506172, 4765.42934217865, 4741.12563204803, 4729.92647341006, 
    4687.20026849259, 4621.4309109743, 4508.13667854925, 4341.3568268946, 
    4177.98478159886, 4005.25872151613, 3906.94146546139, 4005.09763382305, 
    4166.76098724753, 4344.88049919357, 4558.74531000079, 4755.74644683015, 
    4900.42546101331, 5020.23355066846, 5077.54360910379, 5120.79031421237, 
    5160.83579239737, 5193.14409415726, 5206.61219451655, 5196.52326319461, 
    5167.22617037761, 5120.97014455396, 5061.33223542536, 4932.60276691009, 
    4737.93184567838, 4543.18313804642, 4394.52300617727, 4120.12534702319, 
    3497.80386638121, 2545.15399661418, 1792.08568572579, 1226.00599959705, 
    383.165427945073, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    2628.78894248753, 3614.03867681088, 3947.9696202806, 4172.71026609992, 
    4065.89147763595, 3886.23132423409, 3687.56110363779, 3693.22697546435, 
    3858.11575872898, 4037.39705917145, 4249.75359059295, 4367.43365084687, 
    4398.669814687, 4447.11564173189, 4460.65127081588, 4477.78594817756, 
    4492.8019031418, 4463.59538304054, 4250.74312183363, 3788.67540146603, 
    3084.39583534452, 2409.66372591208, 2023.11699781815, 1935.05359591651, 
    1296.63473143658, -0, -0, -0, 0,
  1773.53087788063, 2846.51838184123, 3269.09962781092, 3538.11727447984, 
    3548.40853933474, 3506.19044969643, 3460.60798960719, 3415.92016374789, 
    3356.57248983197, 3247.10103852144, 2951.54335844645, 2455.47202655163, 
    1822.02749545516, 1995.7037959589, 2049.5288349498, 1845.28581193715, 
    1197.59005868694, 597.065028833034, -0, 60, 60, 60, 50, 40, -0, -0, -0, 
    -0, 463.933091178488, 1086.87921984415, 1877.46603275016, 
    2579.04349343873, 2696.58866971183, 2696.58866971183, 2087.89843681754, 
    1768.74629726939, 1665.83606808963, 1260.26187003645, 955.482093541401, 
    -0, 100, 100, 100, -0, 0, 2387.05420861712, 4646.45006003548, 
    5378.97619067688, 5500, 5500, 5500, 5500, 5500, 5131.42164293969, 
    4408.87707887845, 4367.22581609495, 4400.79087979414, 4265.72698845849, 
    4001.65156057947, 3873.74738059611, 3724.65249121604, 4074.11008822629, 
    4341.72864660728, 4341.72864660728, 4335.71155723045, 4350.66838495524, 
    4490.20093095558, 4458.68926564114, 4614.87741266078, 4966.97925698187, 
    5156.18860219666, 5319.60771145571, 5425.41328236041, 5485.29658005964, 
    5488.51980281191, 5431.09287643138, 5270.30067467471, 5293.70837986577, 
    5185.68337939675, 4929.93505361582, 4344.53404537921, 4229.58612758544, 
    4137.87792643411, 4375.04240659872, 4399.8354620457, 4230.4138082762, 
    3925.13659581978, 3897.7381659481, 3912.63797247563, 3659.87962070414, 
    4081.19776594979, 4559.1094926979, 4949.8220616601, 5270.68232144922, 
    5397.15684607523, 5415.11030076877, 5453.09537015411, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5387.54933805921, 
    5129.77760708091, 4900.87238900399, 4782.60637270547, 4898.02142218998, 
    4779.07571895829, 4719.60516006837, 4458.67665853922, 4534.40600022703, 
    4599.81193166093, 4730.05794899007, 4858.46398100632, 4908.29712351049, 
    4834.71450955473, 4973.27537294693, 5090.09770600362, 5164.59078869435, 
    5186.36006982689, 5173.60394054019, 5162.98848989196, 5166.07899658481, 
    5155.33432143901, 5168.05146904188, 5197.04859160492, 5212.72843878887, 
    5240.56920586789, 5220.92198690978, 5195.7388573272, 5166.05192112375, 
    5122.06835617179, 5066.42147337406, 5024.03772775666, 4968.88897898168, 
    4936.50491058438, 4914.8887856215, 4889.3051002686, 4890.18492081819, 
    4881.7440500111, 4883.48075995224, 4893.80326753743, 4900.12080858936, 
    4906.80626323672, 4853.20048230267, 4789.72378022283, 4727.75070560451, 
    4694.99049387114, 4661.31390233341, 4628.41236372707, 4578.90534643126, 
    4529.63890147396, 4462.22790007741, 4394.93017370104, 4321.61452622413, 
    4270.57475305538, 4226.54465246402, 4173.49886063555, 4115.4977594387, 
    4044.56056699724, 3966.11148766767, 3894.23001015397, 3800.00282053956, 
    3692.74997916494, 3578.25024288285, 3492.28622605613, 3509.25278625536, 
    3473.03695811381, 3389.70524479563, 3271.21863448484, 3161.32764218368, 
    3152.60307812715, 3247.64262122515, 3376.17978770714, 3530.70087447633, 
    3683.88769846272, 3830.86658433611, 3905.9704656726, 3928.29976237418, 
    3912.30255640299, 3855.76683690324, 3795.1675298633, 3748.53874276015, 
    3709.37148875504, 3611.01796430157, 3400.02812477454, 3085.41840290381, 
    2868.8023047782, 2432.98344617392, -0, -0, 0, 1672.60653893472, 
    2139.41765910293, 2446.52708029563, 2588.66421886065, 2527.56604773732, 
    2569.49952119183, 2370.34756657681, 907.619598094968, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 254.595707418922, 254.595707418922, -0, -0, -0, 
    637.728619557105, 1405.62049400284, 2154.99077098548, 2989.00500657045, 
    3556.31337329979, 3903.31634935985, 4166.62218585917, 4419.18185522252, 
    4646.07928958404, 4807.48302744292, 4873.18260417047, 4845.89116384828, 
    4803.10769897739, 4750.37349979174, 4657.9831226639, 4530.5564593622, 
    4356.73339463749, 4219.87201212516, 4111.25741610017, 3998.72835671082, 
    4013.74894355475, 4185.37256344044, 4392.57432781064, 4628.42202706312, 
    4832.05186446751, 5008.57278401875, 5129.34608545674, 5222.53673010918, 
    5282.54371227006, 5315.27837448514, 5341.99661362393, 5392.47337503814, 
    5338.06330472028, 5283.14521392043, 5245.44109740679, 5200.29605280601, 
    5105.9, 5073.41037318537, 4918.25181896875, 4792.52992255481, 
    4597.87090036017, 4159.92971588937, 3396.05796032939, 2191.85384798669, 
    1323.95643241201, 789.323136480968, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 2110.2736220506, 3053.99500812493, 3520.08166113863, 
    3838.79121048764, 3866.52940667976, 3849.96778678164, 3739.80805783429, 
    3693.22697546435, 4017.07182162825, 4196.26032382139, 4334.99609061486, 
    4382.37905349296, 4399.8823261736, 4398.669814687, 4399.90381946431, 
    4406.46888969258, 4406.46888969258, 4394.04575603827, 4158.52395516079, 
    3624.86334554243, 2843.70732167682, 2224.39217456823, 1836.64791862072, 
    1724.73049891747, 1296.63473143658, -0, -0, -0, -0,
  2019.7, 2903.2, 3261.6, 3498.3, 3482.1, 3434.6, 3387.2978515625, 3343, 
    3290.4, 3190, 2891.2, 2416.7, 1729.7, 1814.1, 1894.6, 1781.7, 1131.1, 
    565.4, 0, -0, 60, 60, 40, -0, -0, -0, -0, -0, -0, 1196.9, 2012.4, 2704.3, 
    3017.2, 3017.2, 2615.2, 2379.1, 2009.8, 1698.4, 1350.5, -0, 100, 100, -0, 
    -0, 0, 2686.6, 4744, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 4653, 
    4549.1, 4557.6, 4457.8, 4201.6, 4027.7, 3930.2, 4249.2, 4568.4, 4652.9, 
    4701.4, 4727.2, 4809.7, 4883.3, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5281, 5500, 5500, 5037.1, 4612, 4337.7, 4222.1, 4358, 4370.4, 4112, 
    3876.2, 3859.6, 4025.4, 3944.7, 4325.9, 4719.7, 5080.8, 5339.8, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5406.9, 5435.1, 
    5500, 5344.9, 5163.8, 5010.2, 4916.9, 4970.7, 4869.3, 4793.8, 4602.2, 
    4696.4, 4779.07568359375, 4925.8, 5019.6, 5031, 5008.7, 5081, 5175.1, 
    5225, 5220.7, 5213.8, 5202.7, 5215, 5223.5, 5233.2, 5248.4, 5255.4, 
    5269.1, 5248.4, 5214, 5172.2, 5108.1, 5043.6, 4998.1, 4949.6, 4923.7, 
    4909.5, 4898.1, 4896.3, 4891.5, 4884.4, 4891.4, 4901.9, 4913.1, 4868.5, 
    4815.8, 4758.7, 4723.4, 4686.7, 4644.4, 4593.3, 4537.8, 4469.6, 4395.4, 
    4323.1, 4264, 4228.5, 4177, 4129.1, 4065.89135742188, 4000.2, 3938.9, 
    3845.6, 3744.3, 3649.8, 3568.4, 3550.6, 3495.3, 3410.3, 3280.2, 3160.6, 
    3136.6, 3222.2, 3342.5, 3483.5, 3632, 3784.4, 3902.5, 3958.1, 3960.3, 
    3922, 3839.4, 3736, 3620.3, 3483.8, 3272.7, 2950.1, 2513.9, 1380, -0, -0, 
    629.357010774005, 1625.4, 2078.4, 2505.3, 2744.3, 2853.8, 2866.4, 2722.9, 
    1875.6, 270.610395222517, -0, -0, -0, -0, -0, -0, 447.336829274228, 
    447.336829274228, 1027.5, 1027.5, 110, 130, 380, 1009.9, 1617.1, 2324.3, 
    3225.8, 3835.5, 4193, 4426.5, 4627.6, 4794.2, 4887.4, 4907.6, 4859.7, 
    4780.9, 4676.2, 4520.2, 4338.1, 4158.4, 4068.7, 4090.3, 4112.2, 4225.9, 
    4419.181640625, 4627.5, 4849.8, 5042.8, 5207.3, 5314.7, 5361.3, 5500, 
    5407.6, 5500, 5500, 5393.9, 5311.1, 5242.1, 5172, 5105.9, 5044.1, 4934.4, 
    4824.2, 4631.7, 4155.2, 3358, 2133.3, 110, 50, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 840, 
    1192.30999269877, 1203.90872084315, -0, -0, -0, -0, 1478.68884277344, 
    2540.3, 3007.5, 3452.3, 3667.9, 3785.6, 3778.6, 3850.4, 4103.2, 4249.3, 
    4335.1, 4351.7, 4346, 4334.7, 4332, 4339.1, 4350.9, 4316.5, 4046.8, 
    3482.6, 2646.9, 2035.5, 1630.3, 1478.68884277344, 110, -0, -0, -0, -0,
  2265.89457779724, 2959.87331716286, 3254.13644939875, 3458.54161016757, 
    3415.8153998385, 3363.06442869477, 3313.77720860968, 3270.05975048674, 
    3224.31176483909, 3132.84312898806, 2830.93092340047, 2377.92273442567, 
    1637.30133969151, 1632.44385604505, 1739.57882126787, 1718.06075328371, 
    1064.68843747167, 533.667254372407, 0, -0, 60, 60, 40, -0, -0, -0, -0, 
    -0, -0, 1306.87338216973, 2147.3500983973, 2741.96648004957, 
    3337.71512248223, 3337.71512248223, 3142.49304737176, 2989.49028738773, 
    2353.83646468145, 2136.60976946541, 1745.61525880648, 190, 140, 100, -0, 
    -0, -0, 2986.18295581832, 4841.51363606355, 5411.22766443812, 5500, 5500, 
    5500, 5500, 5500, 5347.05920824198, 4897.21976911227, 4730.9498628802, 
    4714.31515339051, 4649.83022140814, 4401.58687980974, 4181.72610745891, 
    4135.82641081598, 4249.2, 4568.4, 4652.9, 5067.16305254663, 
    5103.79050925837, 5129.18954604513, 5307.95501707708, 5456.19024675478, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5291.68685882224, 
    5427.08457411232, 5335.78712274284, 5144.35292642091, 4879.4862726575, 
    4445.82032179472, 4306.40279436646, 4340.97873692566, 4340.97873692566, 
    3993.68341076035, 3827.24395406867, 3821.53384733546, 4138.19383485143, 
    4229.53141738629, 4570.64825060773, 4880.37457734192, 5211.72254648548, 
    5408.95235573718, 5465.3398796307, 5469.41589455698, 5498.55886886849, 
    5500, 5500, 5500, 5500, 5489.60810808337, 5300.98953767046, 
    5279.2626371631, 5313.74513696254, 5370.19934637564, 5396.44759921943, 
    5302.19269689209, 5197.7736435258, 5119.51560720456, 5051.21526989788, 
    5043.30884646315, 4959.46165441282, 4868.06407060988, 4745.64572853883, 
    4858.39838573243, 4956.27846811124, 5121.49888559227, 5180.82233363487, 
    5153.61647783873, 5182.59176454201, 5188.78898213551, 5260.16786141503, 
    5285.50773250036, 5255.01067226852, 5253.96639137917, 5242.45121006526, 
    5264.01633565859, 5291.60964539315, 5298.34860552014, 5299.66867532314, 
    5298.0457367948, 5297.6659466662, 5275.91743201798, 5232.29017176544, 
    5178.31130384232, 5094.12201871462, 5020.79865206129, 4972.08002153156, 
    4930.25072045826, 4910.97440778035, 4904.17070434917, 4906.95444514551, 
    4902.37812734924, 4901.28749179424, 4885.22705941953, 4888.91696537036, 
    4903.77189060196, 4919.40731553427, 4883.72664216888, 4841.8291158718, 
    4789.73462957355, 4751.79600733049, 4712.15879527372, 4660.45066043001, 
    4607.70285941367, 4545.86109546537, 4476.96699500719, 4395.93615834196, 
    4324.6774960402, 4257.45676580896, 4230.43504736873, 4180.51867562791, 
    4142.66727523643, 4086.00247208646, 4034.20248637051, 3983.62971075811, 
    3891.22404341287, 3795.81480508427, 3721.27612304688, 3644.5684130617, 
    3591.86691801513, 3517.57128211319, 3430.80841365764, 3289.09264785582, 
    3159.82850660192, 3120.62482610527, 3196.75856231686, 3308.80106754242, 
    3436.38970720694, 3580.03599777253, 3737.99328373275, 3899.04518960637, 
    3987.981072628, 4008.2840597783, 3988.26007509205, 3883.70768709676, 
    3723.51730899739, 3531.31617697446, 3356.56842942938, 3145.4125718165, 
    2814.71509805255, 2159.06564546907, 326.990295410156, -0, -0, 
    629.357010774005, 1578.15905966602, 2017.3839837057, 2563.99597154131, 
    2899.94680901609, 3180.10165280274, 3163.23403385716, 3075.46605823547, 
    2843.59302194875, 2433.65767814173, 1909.45078312811, -0, 
    1141.25424119393, 1135.67207557004, -0, 1889.19531325076, 
    2265.08606276229, 2252.55712357694, 2212.89581036104, 1800.39886943706, 
    1440.22304006484, 1267.32460139448, 683.282409667969, 1382.06538889809, 
    1828.6277912429, 2493.68308457345, 3462.62822389292, 4114.65164022678, 
    4482.60992261073, 4686.29318862618, 4835.97524545208, 4942.24704475812, 
    4967.39338793996, 4942.07253074219, 4873.45125642641, 4758.61813748609, 
    4601.94742176187, 4382.42429006895, 4145.72677945792, 3960.14985976233, 
    3917.50563412648, 4069.25820603062, 4225.69035100224, 4438.0884476229, 
    4644.90710567176, 4862.44378449506, 5071.12647507689, 5253.53700557306, 
    5406.12425841537, 5500, 5500, 5500, 5500, 5500, 5500, 5449.70796289607, 
    5339.04889415898, 5238.7432005795, 5143.62276148705, 5068.36874964226, 
    5014.87074218205, 4950.57070563957, 4855.86452563469, 4665.60371148298, 
    4150.54559007974, 3319.87548941815, 2074.72373142883, 110, 50, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 466.660196631604, 840, 1320, 1520, 1740, 1740, 1503.6456070567, 
    -0, 840, 2026.70417751144, 2494.90433776173, 3065.78548661781, 
    3469.30002200751, 3721.27612304688, 3817.48484203412, 4007.55904614471, 
    4189.36144784395, 4302.31566430524, 4335.22979127195, 4320.93911197574, 
    4292.09924859968, 4270.77628559023, 4264.12260158398, 4271.65480448291, 
    4295.34868663542, 4238.92910500624, 3935.16868383413, 3340.30801654423, 
    2450.10774805292, 1846.55331367388, 1424.00854822416, 1218.85006590639, 
    110, -0, -0, -0, -0,
  2191.85384798669, 2995.36034946065, 3230.61582387771, 3347.83655593333, 
    3347.83655593333, 3290.34907275594, 3236.89468003951, 3189.34667043156, 
    3144.08042348548, 3077.94212145954, 2770.07458417241, 2371.15996913427, 
    1604.60189521118, 1546.93420037499, 1438.00749801852, 1438.00749801852, 
    1064.68843747167, 533.667254372407, -0, -0, 50, 50, -0, -0, -0, -0, -0, 
    -0, -0, 1280.12060546875, 2141.02788988044, 2741.96648004957, 
    3337.71512248223, 3662.07864033442, 3646.19537599709, 3499.23947967877, 
    3124.25384014213, 2846.3489396192, 2245.06839565153, 1612.13811193514, 
    140, 100, 100, 0, -0, 3502.03458158631, 4879.77500718481, 
    5353.30951773157, 5500, 5500, 5500, 5500, 5500, 5329.18782820277, 
    4828.02122478078, 4796.95550277735, 4821.39086127432, 4748.37091257801, 
    4555.2562480095, 4325.27077971927, 4225.30465018287, 4155.58230441502, 
    4232.53951332936, 4383.89993270823, 4822.96321470744, 5103.79050925837, 
    5343.75447620671, 5343.13497811819, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5364.40096205356, 5488.76870039134, 5331.60931281259, 
    5165.88105371686, 5036.11549112535, 4726.48478950825, 4646.62182990307, 
    4632.5528482721, 4444.9218034671, 4330.18358502389, 4191.11739405576, 
    4294.88396230265, 4383.69557543413, 4528.08824825054, 4825.5127293435, 
    5082.73570232471, 5342.94459911015, 5438.61113384997, 5449.09043028673, 
    5402.21362394666, 5421.78351751197, 5500, 5500, 5500, 5494.72635634689, 
    5350.31404713349, 5088.20127478347, 5126.9783348302, 5253.86031717489, 
    5349.62354864503, 5365.1593951742, 5329.75835088412, 5296.9878079777, 
    5228.72359617158, 5193.92466801967, 5112.79290088618, 5003.92353265576, 
    4943.17197770143, 4945.98623781941, 5056.88531167425, 5170.72935473731, 
    5282.15615908006, 5320.94518446651, 5320.78501289748, 5305.50275830658, 
    5279.98808913006, 5357.59331461891, 5360.1200270531, 5310.97638161736, 
    5317.21200897571, 5336.18716663513, 5357.88751180648, 5372.66093584863, 
    5352.86002495807, 5329.15791694302, 5322.34190790936, 5313.27406593085, 
    5288.22693305497, 5233.2412171454, 5170.96116424993, 5088.6746772776, 
    5020.56339081222, 4934.11432450967, 4914.46807594974, 4905.44175264819, 
    4896.59267742048, 4893.90277890422, 4895.12416076619, 4880.52245950223, 
    4867.13105640703, 4885.0013647046, 4916.2319004955, 4930.72103409461, 
    4911.79152563104, 4851.71289646114, 4797.35721146357, 4753.30297330364, 
    4717.86638462074, 4660.29903486677, 4604.96000237887, 4535.87525005128, 
    4463.72228134859, 4377.17633757161, 4297.12743009457, 4240.59670404025, 
    4205.35943184636, 4171.21785173973, 4130.45627014707, 4094.1632717097, 
    4046.62186928269, 3999.81460710258, 3917.16599867563, 3830.45473934453, 
    3724.53762094, 3691.77812292609, 3644.67368072827, 3571.26425681485, 
    3452.70709436116, 3298.16463478607, 3163.46133715469, 3118.24693977525, 
    3186.05625353942, 3293.11173601181, 3406.16651884114, 3516.75405021977, 
    3655.07227258947, 3826.55783225851, 3960.31826722632, 4036.594649746, 
    3939.77250844097, 3758.79055749512, 3602.7127942859, 3455.03708090591, 
    3292.05602712599, 2777.20382577651, 2106.30119340294, 1520.46475695274, 
    -0, -0, -0, 315, 1130.50552389005, 1697.12502302956, 2401.93688254015, 
    2889.61470802977, 3213.17348883857, 3388.14139621574, 3387.2978515625, 
    3296.04901768248, 3070.86325861669, 2520.38946533586, 1911.17837040794, 
    1642.26087000498, 1628.82052886222, 2077.89636285058, 2599.60312651654, 
    3010.57590635005, 3019.82335640513, 3019.82335640513, 2496.20202873233, 
    1900.80687727448, 1825.89600644411, 930, 1743.98529378248, 
    2047.62106067698, 2693.74915153634, 3672.72668525242, 4286.80425921401, 
    4662.68449464053, 4849.04323227647, 4946.32800024989, 4999.99979033349, 
    4994.76923763902, 4923.36373948309, 4793.817584129, 4648.80885655441, 
    4439.84547982795, 4186.96877121671, 3941.50531787577, 3779.29661939006, 
    3881.01007592347, 4127.37504958626, 4382.4704669919, 4619.96885929813, 
    4843.64377262714, 5066.34422529865, 5260.32465948441, 5434.74985999868, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5428.85883416836, 
    5298.53597925901, 5159.56169536475, 5023.59217787326, 4913.96293658895, 
    4847.57253664582, 4837.94934954173, 4779.07571895829, 4609.89203645817, 
    4089.34774853934, 3282.83927316433, 1968.22781420808, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 466.660196631604, 840, 1320, 1520, 1740, 1975, 1975, 1975, 
    1637.11666950864, 1907.51591205259, 2120.13749152705, 2640.14569793096, 
    3315.54531823347, 3606.25932325728, 3764.36415657999, 4043.8584018707, 
    4201.97327038975, 4278.84568362047, 4298.43406151962, 4261.74791027573, 
    4222.46500851031, 4196.66178003313, 4190.36717320374, 4196.94084824513, 
    4216.92077747017, 4145.17420433891, 3838.55293187736, 3210.37607912572, 
    2311.62757849276, 1737.43435879323, 1424.00854822416, 919.588066567606, 
    -0, -0, -0, -0, -0,
  1645.94981185948, 3052.6495112384, 3234.3821999214, 3334.06268100284, 
    3269.71433372539, 3225.30259771648, 3159.35750915897, 3108.47953191334, 
    3067.89632458945, 2996.08954264528, 2792.52834364938, 2379.02761607198, 
    1343.36035346787, 1343.36035346787, 1306.92062591585, 1436.65273358667, 
    779.752055845596, 350.506003246512, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 924.693080469227, 2029.22779157189, 2578.36642677146, 
    3312.62048461689, 3646.19537599709, 3918.63611177246, 3893.93445065511, 
    3678.08371508891, 3412.36225651085, 2824.82923088048, 2334.8391579467, 
    190, 100, 100, 0, 2013.41442402149, 4399.925713488, 4978.02360446494, 
    5337.38653953987, 5500, 5500, 5500, 5500, 5500, 5346.42515595878, 
    4601.14468817482, 4813.1912838381, 4883.8962757194, 4784.89022555938, 
    4657.81916076801, 4457.70275630036, 4398.75523792748, 4026.37299066266, 
    3874.93739966591, 3903.75541363437, 3660.81342498328, 4966.45432203002, 
    5500, 5271.52056403669, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5331.78153112777, 5500, 5447.7342109732, 5385.39788085709, 
    5214.82369830447, 4861.33399550804, 4730.21179105899, 4640.85717214649, 
    4457.2484779721, 4640.7054783684, 4590.1429086567, 4633.48625946352, 
    4729.39647352861, 4729.39647352861, 5116.37242390443, 5254.9632755972, 
    5427.36453241462, 5500, 5435.14161630998, 5011.52847698748, 
    5279.28000567471, 5469.31274493537, 5500, 5500, 5481.88994650131, 
    5209.59512221045, 4959.73179681908, 5065.85438818348, 5252.26821803902, 
    5224.96594723803, 5408.68565299872, 5436.3826134543, 5407.64230146045, 
    5365.71119180227, 5320.84477027939, 5112.79290088618, 5014.03897425481, 
    4986.01984866688, 4863.18737268082, 5228.56411897088, 5312.91467978129, 
    5437.4861722479, 5446.24159331535, 5453.22903866718, 5390.95907217983, 
    5376.78260524809, 5448.08538727294, 5348.59388653828, 5394.43706941796, 
    5400.69650643197, 5434.62533994295, 5470.87445757078, 5485.69182473469, 
    5380.03836576903, 5371.18168688075, 5347.16946849392, 5325.70839292074, 
    5307.6300504989, 5240.54138874779, 5159.09251766886, 5071.60996988563, 
    5026.97570074346, 4937.20442969887, 4922.2047196466, 4887.5413615739, 
    4873.5960602566, 4857.74451457494, 4841.82303982898, 4835.44865376652, 
    4845.52949100143, 4888.42325104962, 4934.39011287994, 4969.15865770075, 
    4949.78354133204, 4849.48843696928, 4797.37622942677, 4749.41129806859, 
    4694.19910713867, 4636.23401371026, 4610.59527717698, 4535.06041885812, 
    4443.42770918556, 4347.84319245934, 4253.12637373401, 4236.43997758363, 
    4165.4604172959, 4164.37958638672, 4133.21072536682, 4081.78067769336, 
    4046.62186928269, 3980.54321584663, 3951.7639044176, 3851.43325566295, 
    3844.78080778336, 3763.0218244108, 3704.52812421648, 3604.6750312023, 
    3471.95690184006, 3297.4429076298, 3144.39408863866, 3080.09084787914, 
    3176.36903865746, 3300.89700778973, 3391.12041651744, 3451.0287576828, 
    3570.11688943936, 3725.28910694006, 3905.367200348, 3914.33562924143, 
    3799.80988221323, 3695.32866539305, 3642.04549035127, 3524.99113146969, 
    2382.85591468817, 1568.95064190398, 1144.13079789626, 812.827241933817, 
    -0, -0, -0, 0, 667.465769848715, 1526.42978552031, 2122.41796946628, 
    2830.62969656123, 3199.86805480504, 3566.8125059599, 3619.59452711094, 
    3596.29562660768, 3504.54168825436, 3065.78548661781, 2509.85030771973, 
    2161.94790619434, 2107.2883568986, 2600.33084965277, 3143.13431136365, 
    3706.71726668993, 3706.71726668993, 3640.68421741847, 2939.29074980137, 
    1982.279364368, 1982.279364368, 1190, 2019.37882115856, 1952.82084266674, 
    2879.41557615031, 4069.33393715699, 4547.33299501925, 4833.04992412118, 
    5022.99632706945, 5037.16313189929, 5044.58783603241, 4972.00295715528, 
    4852.00945023461, 4688.72802797764, 4524.79325762529, 4261.3301556577, 
    3998.3132615486, 3723.88139113395, 3559.27337916343, 3884.28192771365, 
    4202.59786925099, 4532.27153467699, 4821.36585630985, 4998.39588005439, 
    5240.92127527421, 5377.31011718286, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5378.40824448279, 5218.90275940705, 5054.32297940856, 
    4843.96845685409, 4692.85531828439, 4624.64555527177, 4603.94158748653, 
    4624.06595214262, 4501.64754938763, 4018.51621640591, 3369.73592182211, 
    1533.30779961554, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 766.98377146606, 
    1371.83995867462, 1683.66943352493, 1975, 2235, 2235, 2525, 2525, 
    2353.77382618281, 2693.19428244389, 3333.35267733601, 3524.79447695383, 
    3635.79477153638, 3962.88935542094, 4185.18650483364, 4248.0980069708, 
    4241.32943476456, 4195.4867311102, 4153.02469181273, 4123.17005853551, 
    4115.70689003646, 4121.52043774014, 4140.26500442626, 4090.40912733358, 
    3844.14488192995, 3133.76225357504, 2121.30429160781, 1500.14888152348, 
    1243.94170789094, 565.785293277648, -0, -0, -0, -0, -0,
  2208.19021850232, 2833.15688730094, 3036.56148469188, 3208.64320290215, 
    3211.2423997288, 3146.32489160453, 3079.43690370321, 3021.10108566029, 
    2972.79183688223, 2913.83121032286, 2705.93509710698, 2379.02761607198, 
    1710.07632338801, 1322.16897471123, 1035.70890166586, 838.404972191926, 
    567.197009878129, 343.182678048642, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 924.693080469227, 1796.89069476085, 2297.26815238269, 
    2758.41088867188, 3460.53250614859, 3786.05944386594, 3854.87882347895, 
    3874.29852782887, 3612.96021686327, 3225.36874229647, 2635.71538603206, 
    190, 0, 0, -0, 2596.56009319561, 4226.35066930927, 4898.47888219193, 
    5317.20258256888, 5500, 5500, 5500, 5500, 5500, 5212.56262709074, 
    4601.14468817482, 4839.2603327002, 4908.14950204606, 4932.8213361855, 
    4813.89176716254, 4615.57884811535, 4436.09595229324, 4188.83532809517, 
    3856.303064223, 3831.82492029479, 3660.81342498328, 4225.22534835465, 
    5159.65578078407, 5383.89759557766, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5469.72972298434, 5480.84985415573, 5473.2631815812, 
    5370.89207008801, 5167.63010139224, 4912.53737878112, 4881.14500344442, 
    4640.85717214649, 4668.27489828673, 4730.41806991114, 4703.34977821493, 
    4595.41182694838, 4902.63774542189, 5059.44073169818, 5250.5428338287, 
    5350.31726311806, 5440.6675169844, 5370.10124279321, 5223.58694354815, 
    4902.2472105972, 5015.63711676824, 5193.28430843839, 5336.63281126429, 
    5422.41239955513, 5342.16944501147, 5221.51893433406, 5108.39334777633, 
    5143.41858983545, 5236.5497699308, 5361.8609746499, 5386.27749449299, 
    5410.68108163004, 5351.6771668451, 5241.23636093442, 5118.9904471637, 
    5072.78127383243, 4966.70632817144, 4958.54097728476, 5030.83828748061, 
    5271.13603173922, 5405.65101350138, 5490.85467189437, 5500, 5500, 
    5499.43301217388, 5500, 5488.40108762592, 5481.47955527372, 
    5474.71031128515, 5477.22397000594, 5500, 5500, 5500, 5426.19999736419, 
    5351.9273907179, 5319.36179741107, 5310.86780954052, 5288.2114610505, 
    5254.95044419538, 5190.9056392923, 5126.14690623293, 5066.3354095741, 
    4995.4673327525, 4939.09756064328, 4893.58345999977, 4854.14379867012, 
    4831.83229991258, 4827.03192750398, 4826.13840445955, 4870.84108006908, 
    4902.99077245457, 4943.79413429631, 4972.72331121348, 4944.03499283915, 
    4873.70350295518, 4794.51390169872, 4726.2687190164, 4663.30832410519, 
    4600.51016187961, 4546.27145541936, 4470.47508169263, 4380.96186801868, 
    4283.10340982093, 4179.68181910339, 4160.57571713161, 4126.29268285838, 
    4107.25175804882, 4079.9564191392, 4038.50394469985, 3989.85211225899, 
    3923.13092131826, 3856.60570939427, 3778.06820151658, 3721.27612304688, 
    3723.66995360483, 3676.39159213909, 3613.69720447034, 3445.72916135273, 
    3287.73537532978, 3166.74533421229, 3159.80333894026, 3241.79565047996, 
    3348.20206408611, 3419.41329078905, 3438.95409878586, 3504.20893182607, 
    3599.61852266999, 3659.67189754352, 3636.13591466105, 3585.28021752949, 
    3407.40665713879, 2964.89675127163, 2362.9933921818, 2119.78450300097, 
    -0, -0, -0, -0, -0, -0, 0, 606.500040516954, 1128.50636549985, 
    1673.93336823849, 2376.23456005716, 2873.44466450477, 3340.48340631071, 
    3599.51211081135, 3649.54873322289, 3537.11807672992, 3366.83589748997, 
    3103.90760523265, 2990.92947593754, 3168.98592294393, 3510.3279261156, 
    3894.51672157795, 4144.08669919501, 4192.04347592029, 3753.83233865981, 
    3170.70385737566, 2377.20020213438, 2178.89011346403, 1190, 
    2162.64690548682, 2669.55655341437, 3407.70215723366, 4245.60375582131, 
    4750.78056339049, 5042.98007243473, 5116.40335947914, 5116.40335947914, 
    5037.5027611662, 4903.98045166623, 4734.6797623333, 4522.71486867552, 
    4291.44366601853, 4027.67620174655, 3809.48228592631, 3629.76880880965, 
    3652.98714419684, 3942.40259349278, 4259.48192236503, 4578.79456120881, 
    4837.75070655764, 5046.00629338344, 5236.92920538434, 5382.80321412541, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5480.57201810854, 
    5315.6246675385, 5123.32958177759, 4883.10619926195, 4615.13003413868, 
    4369.2428475504, 4270.91893685978, 4267.47622829531, 4301.65722205383, 
    4218.96084654172, 3729.62905927495, 3083.72004931323, 1533.30779961554, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 1458.24515816833, 
    1548.04978716056, 2235, 2235, 2525, 2525, 2525, 2693.19428244389, 
    3038.42810398504, 3311.81307646858, 3571.50109040824, 3847.48835701732, 
    4048.09260122729, 4150.96700207967, 4143.27270554989, 4098.07662784766, 
    4075.06652803667, 4045.20559928236, 4035.72135211953, 4040.80252949303, 
    4048.70595669214, 3959.79356132966, 3654.54288399168, 3018.50096187769, 
    2121.30429160781, 1610.50925363485, 1044.89927061619, 565.785293277648, 
    -0, -0, -0, -0, -0,
  1862.58654731823, 2763.48806395647, 2949.14676948003, 3065.78548661781, 
    3135.56784859283, 3065.78548661781, 2986.79648890033, 2923.04066114943, 
    2882.58818419774, 2814.39884551037, 2692.18933375695, 2439.88392868226, 
    2062.71189963643, 1051.47380257324, 654.612458198456, 441.792810096934, 
    308.468064719436, 190, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    722.69558750426, 1367.50588413406, 1948.80465477325, 2508.2158671771, 
    3108.78141632672, 3793.80532646816, 3907.02097301736, 4034.45672090155, 
    3899.50434049713, 3627.34761400679, 2762.76304809381, -0, -0, 
    1007.94216597725, 1657.54963760261, 3035.17259889014, 4326.8558534928, 
    4960.75985711723, 5322.72872895582, 5500, 5500, 5500, 5500, 5500, 
    5120.08621519413, 4588.00982882201, 4848.14894624072, 4949.84909166527, 
    4894.74539267209, 4829.79076514482, 4752.88774809199, 4623.21306059717, 
    4354.84601469421, 3698.95956548843, 3599.31982456083, 3609.54840717973, 
    3387.2978515625, 4665.71481152995, 5500, 5480.86583058826, 5500, 5500, 
    5500, 5500, 5500, 5489.15812678147, 5500, 5385.10720267987, 5500, 5500, 
    5401.99665027083, 4993.78509593915, 5088.87456443707, 4985.37687128531, 
    4800.76252425272, 4958.35863559203, 4765.29047276236, 4942.40460262666, 
    4930.85937415241, 5072.99589926845, 5097.5358928567, 5408.86324369995, 
    5451.81359048847, 5443.60391337401, 5357.26587883543, 4956.97144329587, 
    4609.2898239409, 4558.18815635484, 4888.08636422044, 5228.42740433769, 
    5235.67037380359, 5363.31363895264, 5315.12369410172, 5111.82177563278, 
    5164.87587947778, 5206.32188755652, 5411.70153619676, 5258.62747936645, 
    5467.61235769298, 5422.61979349681, 5227.25829028908, 4928.53327300269, 
    4884.48304451863, 4947.89335760516, 4918.03789632009, 5196.42124379521, 
    5385.92922586452, 5493.32964530684, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5476.24299578138, 5500, 5500, 5500, 5447.2479064153, 
    5318.88120831885, 5308.14443453066, 5369.60741732193, 5282.20204053541, 
    5272.28302561599, 5209.83552428512, 5132.11934070115, 5110.82038752857, 
    5034.17765668431, 4976.60584355559, 4910.64281700449, 4863.64314349401, 
    4847.87706026031, 4832.73085349134, 4872.58628067323, 4888.3112926103, 
    4906.64244631634, 4967.15125724518, 5011.45873671296, 4961.64057371957, 
    4877.16928297713, 4779.07571895829, 4693.9681471866, 4608.26064946132, 
    4552.97889428238, 4469.85298134419, 4419.18185522252, 4357.55676718331, 
    4250.63772498847, 4173.56189720487, 4142.38297601575, 4092.34592504642, 
    4070.80125500474, 4041.21925066322, 3983.39819443791, 3936.70231670377, 
    3848.92960333278, 3780.63433607516, 3660.86988045223, 3531.53566361877, 
    3676.39159213909, 3703.11748927293, 3592.31529281117, 3436.46233422929, 
    3271.72803872694, 3131.02565093345, 3191.33858918372, 3324.709834762, 
    3359.1269092785, 3395.6772589238, 3402.22592420559, 3375.86473384553, 
    3449.34655495723, 3534.27039959755, 3578.18458918748, 3578.18458918748, 
    2320.34746833347, 1559.11602584742, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    334.000057365342, 1575, 1575, 2111.67413344319, 2371.02272402902, 
    2858.50730952754, 3553.94351880276, 3553.94351880276, 3537.11807672992, 
    3392.07443671563, 3387.2978515625, 3456.32201162042, 3721.27612304688, 
    4033.52264621214, 4347.5242324891, 4626.45897627842, 4593.41113923563, 
    4049.12966509738, 3273.03818025372, 2264.24661185372, 2315.20251902575, 
    1190, 2346.25893103586, 3175.60391349151, 3784.31338351774, 
    4759.77671955393, 5097.88088936825, 5263.82823717944, 5280.94508423178, 
    5172.01856245335, 5045.19063359983, 4823.05334892292, 4655.64920464047, 
    4382.95031187079, 4022.33489074374, 3836.43046475282, 3647.70822344409, 
    3470.07086632297, 3615.04688800488, 3986.14146126372, 4338.24326728985, 
    4670.76397256519, 4890.77732921888, 5047.99020885445, 5275.41472404896, 
    5452.16470644575, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5435.08832744298, 5231.87914203399, 5042.18104975027, 4731.55517453957, 
    4352.586865846, 3840.94675696527, 3835.01582541905, 3955.17811208586, 
    4023.36342728658, 4023.36342728658, 3598.1954230288, 2924.56953535332, 
    1511.92347607909, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 280, 280, -0, -0, -0, -0, -0, -0, 
    1304.01344512848, 1774.32243192946, 2525, 2525, 2525, 2589.64582115205, 
    2842.07092517115, 3128.36523512269, 3507.15082004857, 3796.85169750991, 
    3990.21981785971, 4092.16477571436, 4070.07255810876, 4032.72087541006, 
    3996.72751052042, 3959.31978942172, 3936.90035793103, 3947.6951462356, 
    3962.23334046544, 3894.47534479396, 3664.10109695471, 2959.17208959572, 
    2118.83222549113, 1638.39507048552, 683.282409667969, -0, -0, -0, -0, -0, -0,
  1727.16632973362, 2333.8583813939, 2647.01499166251, 2859.85950887346, 
    2923.78398536632, 2957.5500696347, 2896.40601178629, 2828.4169561149, 
    2772.46753788719, 2711.76885842095, 2624.20474123011, 2384.29334313699, 
    2015.40255384164, 1328.74737794075, 765.839862443459, 436.718704624532, 
    253.361404418945, 150, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    706.54528222211, 1087.18481613606, 1547.08767414927, 2191.85586547772, 
    2794.13183215302, 3322.4816767568, 3791.13679976805, 3884.64813940851, 
    3808.40942217885, 3563.11481522854, 2925.90431624904, -0, -0, 
    2084.48894936648, 2665.05368962119, 3547.54183009883, 4326.8558534928, 
    4887.90795584822, 5251.64131745859, 5432.23002765998, 5500, 5500, 5500, 
    5434.31822373961, 5120.63557617372, 4796.43063328634, 4856.40292714631, 
    4902.39419243567, 4931.40053070079, 4863.15274845805, 4779.07571895829, 
    4600.40604803427, 4298.33538688301, 3864.43297664329, 3489.73607834033, 
    3496.00908118914, 3502.66664684497, 4322.7957811565, 5048.55254313621, 
    5212.19448832136, 5438.93168534732, 5500, 5500, 5500, 5500, 
    5411.70944878543, 5463.3637900179, 5500, 5500, 5500, 5339.18764217477, 
    5033.44967848779, 5089.68673221586, 4975.24426069192, 4890.57935216777, 
    4970.2167719406, 4945.23367149194, 5007.13906083144, 5148.8429516224, 
    5171.70856508181, 5249.9950902667, 5342.52547444766, 5350.70847053786, 
    5277.96290417772, 5174.00015208862, 4935.51688145589, 4644.94758468016, 
    4509.41855984438, 4654.1434824032, 4957.69998567515, 5168.04355130616, 
    5205.4658779784, 5148.13019600496, 5019.83962925825, 5093.6122585064, 
    5189.91839934915, 5256.90486391223, 5308.53779299965, 5305.78961057284, 
    5143.41858983545, 5028.5229974399, 4885.29757451611, 4825.4116090142, 
    4874.60384782916, 4968.79110633712, 5215.4551642048, 5369.67600049009, 
    5472.38905382749, 5500, 5500, 5500, 5500, 5500, 5447.24437685293, 
    5392.45512947336, 5391.54651353238, 5424.07590906773, 5493.37171261711, 
    5500, 5495.84924389989, 5426.05924763055, 5351.51097331798, 
    5338.71054599251, 5325.84088831705, 5319.69708656632, 5320.59011126936, 
    5326.44510806228, 5292.55423649965, 5243.60085891672, 5155.87662673792, 
    5085.62479152425, 5009.27845468254, 4958.58377599629, 4928.58760755921, 
    4914.38997623062, 4902.43460685823, 4894.31184936761, 4936.43581688517, 
    4972.61304667558, 4986.88544429828, 4953.94265379911, 4888.46647932993, 
    4797.82850331146, 4700.29968195082, 4592.69329954737, 4512.48208441492, 
    4428.37666316664, 4362.01932885618, 4269.02594179929, 4185.74307108585, 
    4107.45482216547, 4065.89147763595, 4017.95233213368, 3998.89536610385, 
    3962.47762468674, 3906.60285146125, 3842.58977053713, 3757.07718505366, 
    3668.49336119555, 3562.25802606518, 3547.47313123047, 3619.99403284372, 
    3644.7793959325, 3580.46736935147, 3398.77082323879, 3241.85186333584, 
    3187.68762447508, 3255.85120653322, 3330.52175070313, 3368.25056135553, 
    3359.1269092785, 3355.27828371537, 3354.09000893637, 3366.83630807506, 
    3305.36635761248, 3110.89446885193, 2517.28330630079, 1968.45205878905, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 985, 1575, 1575, 
    1740.36213296567, 2155.96669831801, 2616.52705419852, 3040.73244705194, 
    3397.02177601297, 3602.6605754927, 3523.46689933944, 3498.80301890542, 
    3637.80951620177, 3827.90484040857, 4033.52264621214, 4379.5775056499, 
    4577.89819621845, 4510.66829459361, 4049.12966509738, 3273.03818025372, 
    2378.93958286078, 2209.8611153986, 930, 2803.48938915152, 
    3619.34249476349, 4258.38468196548, 4891.40865906916, 5209.60576488264, 
    5337.86577900889, 5324.8082925678, 5220.06511040104, 5026.2543360696, 
    4779.07571895829, 4419.18185522252, 4105.92657123972, 3895.70334122363, 
    3741.55762539207, 3630.70484026352, 3635.04345289023, 3828.81804676436, 
    4126.27473256786, 4441.56842383448, 4708.27074291839, 4934.54577779048, 
    5092.57082675903, 5206.78194043791, 5305.83377920571, 5387.15511055436, 
    5500, 5500, 5500, 5500, 5496.48793787393, 5397.78007340532, 
    5273.24638792482, 5113.04703290636, 4883.32510154416, 4528.99438024736, 
    4099.06394290306, 3511.56461028608, 3269.01926583604, 3517.22877708608, 
    3762.18774366849, 3756.45298256839, 3424.72222239125, 2824.62653835006, 
    1947.03102490917, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 440, 440, 440, -0, -0, -0, -0, -0, -0, -0, 
    -0, 1705.33803602083, 2092.99425020388, 2320.83130065214, 
    2574.44011974494, 2840.59121082453, 3121.40799210248, 3464.07223247569, 
    3700.50974551931, 3866.10016734519, 3945.669679493, 3974.97931651584, 
    3962.6121655387, 3920.43382972245, 3881.03199721309, 3850.74266385693, 
    3850.2839262796, 3844.48022621793, 3756.91161947502, 3458.94403617891, 
    2873.1003426285, 2121.15361777088, 1478.68884277344, 683.282409667969, 
    -0, -0, -0, -0, -0, -0,
  -0, 1531.05668302307, 2211.44063868916, 2685.11641094177, 2760.08813618268, 
    2780.5914925103, 2768.14148447285, 2706.33719511788, 2651.83619374201, 
    2581.83742295391, 2527.46674242718, 2389.02611180822, 2122.2693935769, 
    1559.46847137778, 683.282409667969, 220, 90, 90, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 311.493373920296, 587.571105970273, 914.338518804828, 
    1173.31789636472, 1700.26313166992, 2466.66776221529, 2576.7950972069, 
    3721.27612304688, 3875.48829053922, 3800.3574897231, 3630.96108464189, 
    2778.48083074288, -0, -0, 2883.93302405136, 3512.71523096648, 
    3516.40613859692, 4115.15581504092, 4803.43197993262, 5025.92977436803, 
    5420.13170477725, 5500, 5500, 5500, 5500, 5352.80206255096, 
    4857.20836619187, 4912.4349336536, 4949.03222515171, 4929.37471198833, 
    4796.25265936816, 4855.81063585565, 4681.98388197612, 4381.17986183252, 
    3897.99519734354, 3452.68681871346, 3425.5998526668, 3295.1130548202, 
    4038.64816830546, 4717.62398833305, 4844.8067282087, 5227.43324885677, 
    5397.63585999683, 5377.79498284148, 5347.87939387254, 5420.60054530274, 
    5369.11910159207, 5173.84357529143, 5500, 5500, 5500, 5500, 
    5291.90806912934, 5225.68489312495, 5075.98120501103, 4982.75923768619, 
    4981.03019806581, 5081.07269397218, 5091.73264708263, 5176.12310950204, 
    5262.12347775747, 5312.64655929565, 5237.6849785946, 5181.64489626365, 
    4867.27447543009, 5034.77713637383, 4812.77751887191, 4419.18185522252, 
    4246.44974690515, 4363.14438898472, 4799.33692597679, 5013.40146276878, 
    5023.26356433575, 4968.60319708117, 4910.06984182582, 4825.87630130442, 
    4986.40472739756, 5009.18006675859, 5163.30069620877, 5271.28405492802, 
    5093.24021901624, 4751.71830452122, 4574.71602499207, 4824.40359309984, 
    4832.11229216962, 5143.41858983545, 5273.53884945193, 5414.42945248425, 
    5471.48158689803, 5470.67128308541, 5433.18703415193, 5500, 5500, 
    5424.94138709317, 5301.46741832732, 5215.35357260674, 5223.59786893631, 
    5290.74702924195, 5391.32981807446, 5440.46694876913, 5420.66926282985, 
    5378.93323872994, 5309.983739699, 5313.62943924043, 5330.64787067363, 
    5336.49656692029, 5379.35773754352, 5388.3617792365, 5373.10834009577, 
    5356.84706887675, 5283.48724917695, 5245.13684255087, 5207.41369491436, 
    5128.73362976064, 5026.31972620823, 4959.82316327152, 4948.4008390415, 
    4911.13660421676, 4961.48250335517, 4973.04142822643, 4996.05542229297, 
    4950.10084337141, 4899.87219495331, 4808.97503808309, 4701.51104522127, 
    4566.00491125984, 4461.21318104134, 4363.09457987885, 4281.80605701901, 
    4155.62301818549, 4103.36042468897, 4013.95702989861, 3990.16764252821, 
    3922.64102862353, 3899.67370563876, 3880.537057547, 3844.10020966943, 
    3741.15711178128, 3654.09056860855, 3545.45519502953, 3343.66593633973, 
    3453.26948802476, 3457.9910821286, 3514.00172397198, 3588.58355488231, 
    3304.75730178413, 3156.34668336859, 3184.2425763965, 3272.19952718472, 
    3336.56759426422, 3359.1269092785, 3359.1269092785, 3355.27828371537, 
    2740.02033354383, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    1386.18433258159, 1455.73514302014, 1455.73514302014, 1227.58171123963, 
    908.121865935783, 1575, 1575, 1575, 1575, 1813.80556903191, 
    2209.32120547588, 2524.16504991724, 2880.37191400961, 3279.08608509058, 
    3367.88384867656, 3367.88384867656, 3677.2883940677, 3825.52894065379, 
    3955.94841000781, 4184.1714964453, 4371.07763156596, 4248.28960300977, 
    3853.04190370226, 3187.73387817806, 2211.44169197477, 2070.63263207092, 
    650, 3235.30484194406, 4259.58505663067, 4901.32318815192, 
    5185.40972525916, 5250.98175392029, 5341.66977822495, 5353.65953636373, 
    5237.44218999206, 5045.47215601393, 4734.29909656036, 4390.80678921734, 
    4114.12620112923, 3900.56817538205, 3635.17967767518, 3472.2036214783, 
    3662.34051615009, 3910.97753316907, 4249.69344064051, 4537.1329107854, 
    4780.70571364158, 4999.1287036622, 5131.95774541632, 5131.95774541632, 
    5099.58254760419, 5173.18733762897, 5284.5345665522, 5385.36249606265, 
    5386.67601627442, 5346.54698014028, 5296.70078052871, 5209.64645522021, 
    5129.83206031607, 4983.81454648242, 4740.70660236295, 4419.18185522252, 
    3975.98737448697, 3531.42050930854, 3218.3863056674, 2880.42490636587, 
    3566.01995092265, 3567.05443003338, 3323.8430338761, 2866.53654734559, 
    2146.59602239835, 1002.87911427475, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 700, 700, 700, 440, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 1748.51366141208, 2243.20434667649, 
    2592.73599623336, 2897.5019880846, 3093.43895273702, 3431.31907466122, 
    3587.41203961898, 3577.60153701829, 3782.8287408313, 3896.77601816852, 
    3887.18377932417, 3833.91207438199, 3783.58305100366, 3738.85194303444, 
    3747.82825038827, 3706.12408977943, 3626.34491361748, 3361.32490811928, 
    2801.22709390739, 1987.4546710214, 1170.74157454671, -0, -0, -0, -0, -0, 
    -0, -0,
  -0, -0, 1796.49617019774, 2272.79175277828, 2511.08596112839, 
    2579.18671183312, 2572.51688947023, 2563.79255434741, 2503.35686900178, 
    2441.34392377011, 2406.03870868304, 2284.66547555935, 2058.74181490373, 
    1559.46847137778, -0, -0, 80, 80, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    255, 311.493373920296, 542.381194560993, 885.466628106794, 
    1131.47462124555, 1554.14654460321, 2295.27346815355, 2626.4, 
    3450.57680774794, 3736.87693045143, 3756.15267434701, 3513.01322517223, 
    2939.29584230155, -0, -0, 2883.93302405136, 3522.90920647022, 
    3559.58362244447, 4266.12517078132, 4741.65270791556, 5098.97901248551, 
    5336.89347372879, 5489.46074442032, 5500, 5500, 5500, 5418.343317597, 
    5108.81315311485, 4961.84023220822, 4911.12824385711, 4894.83802858537, 
    4833.94352081394, 4779.07571895829, 4633.38276205591, 4346.3376425884, 
    3912.70704259323, 3484.71561107517, 3397.83040307056, 3295.1130548202, 
    3873.98941431029, 4676.15998841151, 5064.36955898866, 5091.54947579128, 
    5037.64967233189, 5089.88916115025, 5096.30211455101, 5218.11917211354, 
    5177.73598649884, 5479.98907124146, 5500, 5500, 5500, 5500, 
    5398.60738733011, 5272.39392455924, 5089.30592983723, 5067.62571602437, 
    5085.23097828762, 5014.67835548103, 5063.80847441309, 5056.09012120513, 
    5120.96923695376, 5120.96923695376, 4990.10016321753, 4813.04263812665, 
    4703.08468261889, 4646.29008462504, 4491.51416969893, 4298.04719910119, 
    4212.16508782068, 4323.59217630024, 4560.80166555321, 4745.21371896419, 
    4825.90583527004, 4791.42356545847, 4662.63835077794, 4612.261776144, 
    4573.60309471199, 4725.33458522641, 4880.84595763961, 4942.64582959807, 
    4902.97612762422, 4751.71830452122, 4599.74168489771, 4694.58492419515, 
    4940.263034927, 5168.27463827783, 5328.76003548471, 5428.7640065288, 
    5467.73748392208, 5444.81608866198, 5478.07845430186, 5457.48966812646, 
    5362.57892377398, 5224.42792032635, 5084.33498710457, 5010.94020429691, 
    5028.07880801274, 5113.10536203246, 5236.78416260816, 5310.09224945805, 
    5337.23699052964, 5346.06939785792, 5332.94210937401, 5336.10128304635, 
    5350.10575144837, 5344.87861228223, 5369.03294453431, 5395.1475709626, 
    5398.42679528625, 5400.74738540788, 5380.42458545383, 5344.2211012809, 
    5287.54984824178, 5224.29865924143, 5170.59632610591, 5117.33302447449, 
    5067.87693076503, 5027.83464046845, 5019.23110821328, 4985.46924699761, 
    4984.98578942821, 4958.75832045614, 4882.0267383597, 4779.07571895829, 
    4656.43749782855, 4524.03568332792, 4408.91910864414, 4310.55218706024, 
    4228.5301889847, 4135.1324721344, 4054.09547297191, 3974.63225814259, 
    3949.02624250758, 3895.80552740388, 3835.44626321526, 3817.26925299163, 
    3767.28140372778, 3671.63178283299, 3560.75655751721, 3446.41654677682, 
    3371.64028551422, 3398.21312243673, 3465.25588673561, 3488.81591018929, 
    3480.9820082358, 3317.85285897734, 3167.25065197066, 3148.40358964349, 
    3235.17816875625, 3339.91157214455, 3255.66844956569, 3046.73796482511, 
    2794.79190638344, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    1678.35749210353, 2598.55573540681, 2483.88729780855, 2265.13737147027, 
    1824.40476197392, 1766, 1766, 1575, 1672.50433735539, 1746.54966525087, 
    1935.98581519077, 2191.85384798669, 2466.66776221529, 2844.04607538409, 
    3208.8738507199, 3315.99491271807, 3363.82908434197, 3631.96923235633, 
    3774.73961288713, 3893.60383461698, 3962.62830562957, 3851.56369938248, 
    3496.16492950219, 2878.72824895521, 930, 930, 2243.19147161703, 
    3858.48852713427, 4621.82372098437, 5118.51000269268, 5341.38660706045, 
    5409.74013131656, 5400.61600368734, 5295.23255288263, 5122.3962618183, 
    4929.58274151225, 4684.60438253891, 4430.12436519292, 4139.8779750757, 
    3871.23071897135, 3657.56903859697, 3538.03036454721, 3675.31458918885, 
    3882.44628316892, 4246.6783773625, 4537.91870962726, 4787.52335655908, 
    4996.86788922052, 5158.71411468602, 5228.14316158989, 5258.18345538889, 
    5254.26726624579, 5270.87116654943, 5257.79778176103, 5242.04694189261, 
    5193.73851080318, 5120.92433002593, 5038.59156416521, 4958.29114093888, 
    4835.96211772116, 4603.8838716044, 4249.6608169495, 3673.76710308798, 
    3232.1550556499, 3178.64414338359, 3141.25485085696, 3390.88711846297, 
    3399.28186160391, 3215.75651883758, 2758.41088867188, 2158.8965469637, 
    1002.87911427475, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 960, 960, 960, 440, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 2042.89458956881, 2231.59003205727, 2577.73857171284, 
    2928.30511899891, 3164.3727041397, 3367.37519537361, 3492.12155410135, 
    3736.08608884253, 3808.61103774219, 3804.77704769164, 3753.63085074716, 
    3685.52307138015, 3631.46200034765, 3612.23021683146, 3543.85953787379, 
    3428.6208641578, 3081.71134144258, 2468.93874465024, 1710.94803481647, 
    989.152946303827, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, 308.546024677228, 2098.7, 2284.2, 2318.6, 2308.3, 2245.9, 
    2199.7, 2155.1, 2057, 1912.7, 1550.3, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 254.2, 255, 255, 713.8, 1016.6, 1404.7, 2001.1, 2626.4, 
    3160.2, 3487.3, 3583.9, 3450.5, 2982.1, 0, -0, 3007.2, 3809.2, 
    4065.89135742188, 4538.9, 4847.6, 5144.1, 5368.1, 5494.7, 5500, 5500, 
    5500, 5500, 5281.9, 5018.9, 4914, 4863.3, 4817.6, 4779.4, 4609.4, 4319.1, 
    3890.1, 3517.4, 3409.5, 3363.9, 3855.2, 4557.9, 4967, 4995.4, 4927.7, 
    4962.1, 5071.1, 5237.9, 5285.5, 5500, 5500, 5500, 5500, 5500, 5500, 5183, 
    5054.4, 5042.1, 5032.1, 4985.3, 4992.4, 4987.9, 5068.2, 5011.2, 4719.3, 
    4384.4, 4319.5, 4275.6, 4192.6, 4107.8, 4106.6, 4163.2, 4380.9, 4563.6, 
    4548.1, 4555.4, 4504.9, 4422.9, 4305, 4334.7, 4462.5, 4642.5, 4627.9, 
    4585.1, 4480.5, 4690.4, 4948, 5173.5, 5335.9, 5402.2, 5500, 5500, 5500, 
    5294.2, 5151.4, 4941.3, 4730.9, 4662.1, 4736.6, 4935.8, 5110.8, 5234.5, 
    5304.3, 5334.4, 5346.7, 5355, 5358.7, 5354.1, 5376.5, 5400.8, 5412, 
    5423.6, 5416.5, 5389.6, 5500, 5273.7, 5215.9, 5173.4, 5143.41845703125, 
    5099.7, 5086.5, 5051.6, 5026.1, 4973, 4889.4, 4779.07568359375, 4658, 
    4521.2, 4380, 4281.6, 4202.3, 4119.4, 4065.89135742188, 3992.5, 3938.4, 
    3885.4, 3828.3, 3784.2, 3724.5, 3602.1, 3512.1, 3400, 3312, 3322.9, 
    3391.8, 3420.9, 3391.9, 3229.6, 3086.2, 3042.1, 3010.79207272935, 
    2444.45497030586, 507.103879968353, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 1678.35749210353, 3097.40445097477, 3336.35524950757, 
    3336.35524950757, 3325.79718520838, 3221.51452826348, 1981.95483728453, 
    1815.208380174, 1514.51265784191, 650.169517082769, 708.374842558267, 
    1233.43430080021, 1233.43430080021, 930, 930, 1101.54602050781, 
    1101.54602050781, 3631.96923235633, 3631.96923235633, 3594.31349649527, 
    3545.68869087508, 3612.47968967251, 1350, 1350, 326.990295410156, 
    495.553629324057, 2243.19147161703, 4421.9, 4963, 5294.5, 5500, 5388.6, 
    5330.7, 5197.3, 5044.3, 4911.4, 4720.2, 4495.3, 4210.7, 3936.9, 3689.4, 
    3527.8, 3636, 3865.5, 4228, 4532.9, 4792, 5009, 5179.3, 5275.8, 5500, 
    5318.5, 5289.5, 5230.7, 5184.2, 5094.3, 5011.7, 4928.8, 4859.6, 4751.6, 
    4553.2, 4253.1, 3824.8, 3494.8, 3387.2978515625, 3311.7, 3356.2, 3356.2, 
    3145.9, 2668.3, 2104.1, 220, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 960, 960, 960, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 599.298033095319, 1369.11438702269, 2501.7, 
    3101.5, 3332.5, 3603.3, 3721.9, 3721.27612304688, 3659.2, 3574.6, 3496.7, 
    3459.2, 3373.2, 3165.2, 2700.7, 1963.1, 1114.8, 70, -0, -0, -0, -0, -0, 
    -0, -0,
  -0, -0, -0, -0, 1686.34992647229, 1989.23060319206, 2064.68356578678, 
    2052.8094083634, 1988.49891264665, 1958.09892593535, 1904.18309941917, 
    1829.41444247737, 1766.64054677782, 1403.55286720158, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 200, 253.361404418945, 253.361404418945, -0, 
    542.075624571914, 901.730690814897, 1255.32558363609, 1706.84673621789, 
    2380.74978511648, 2869.77478739174, 3237.78729776682, 3411.67825503374, 
    3387.93298954673, 3024.87799954859, 1650, 2477.89897827202, 
    3130.46832411235, 4095.5342238335, 4572.10397707792, 4811.71186100954, 
    4953.52959651934, 5189.28672921158, 5399.25545462813, 5500, 5500, 5500, 
    5500, 5500, 5454.95361715278, 5075.98913334785, 4916.92133666221, 
    4831.84737929988, 4801.20908777431, 4779.62957399755, 4585.43117215182, 
    4291.9455172855, 3867.47503052471, 3550.11153463094, 3421.26915480389, 
    3432.78312626893, 3836.32398220187, 4439.60409741195, 4869.62520980074, 
    4899.29058539125, 4817.71288130861, 4834.41049114518, 5045.87556478569, 
    5257.7432794244, 5393.31258380124, 5436.3953142009, 5500, 5500, 5500, 
    5422.6942192, 5278.27674486227, 5093.6589116521, 5019.46008667013, 
    5016.5291345804, 4979.01468551512, 4955.98156322132, 4920.90978270601, 
    4919.66354512091, 5015.38519654437, 4901.52742429044, 4448.51528032165, 
    3955.78346362451, 3935.87247391361, 3904.98225695271, 3893.7293122045, 
    3917.5008339296, 4001.05589701596, 4002.79827184394, 4201.04419635632, 
    4382.06723943616, 4270.38244333388, 4319.45520724339, 4347.19006057727, 
    4233.45975220075, 4036.47130717096, 3944.06438634025, 4044.13435105578, 
    4342.27130125645, 4352.83047626022, 4361.20853370258, 4361.20853370258, 
    4686.17653687276, 4955.80435388181, 5178.6641222485, 5343.03333791461, 
    5375.70703681178, 5366.36041131237, 5329.30549022399, 5264.61267963558, 
    5130.92862009142, 4940.20112395139, 4658.20928832995, 4377.56073408715, 
    4313.17036079669, 4445.03918956934, 4758.39851805082, 4984.72211852717, 
    5158.95059289007, 5271.41337526397, 5322.79091189051, 5360.51656680311, 
    5373.82672401071, 5367.22189218261, 5363.27399662938, 5383.98003578549, 
    5406.39380483639, 5425.57293567518, 5446.55003124467, 5452.49580066727, 
    5435.0611819907, 5402.26352231707, 5323.11883918363, 5261.23572945885, 
    5229.4751677329, 5204.09107223181, 5171.58490210823, 5153.78078157979, 
    5117.78620819975, 5067.3095274941, 4987.16640737746, 4896.72522672439, 
    4764.1635758297, 4659.49063060312, 4518.39993283815, 4351.17196279054, 
    4252.58438061632, 4176.1547338788, 4103.65048308682, 4065.89147763595, 
    4010.28998569163, 3927.79202159447, 3874.96618650408, 3821.23914346924, 
    3751.06046002062, 3681.67651642835, 3532.66833360139, 3463.34965430319, 
    3353.55394945165, 3252.38255640819, 3247.65930151504, 3318.28246331373, 
    3352.92545896372, 3302.86247332315, 3141.27040209627, 3005.08543244636, 
    2935.73746145071, -0, -0, -0, -0, -0, -0, -0, -0, -0, 617.3497625183, 
    617.3497625183, 371.797854437214, 0, -0, -0, -0, 1678.35749210353, 
    3097.40445097477, 3336.35524950757, 3336.35524950757, 3325.79718520838, 
    3272.3308995302, 3088.96157275255, 3027.82192117386, 2758.41088867188, 
    2409.66088288634, 2139.56463702486, 1900, 1900, 1492, 930, -0, -0, -0, 
    1350, 1350, 1350, 0, 3258.87780591381, 3083.54545711376, 
    3052.86329944703, 3469.49103263054, 4299.53187626364, 4985.23866196083, 
    5304.10514269152, 5470.40595204751, 5435.75230205482, 5367.46219673319, 
    5260.70129228974, 5099.39485061571, 4966.17359371578, 4893.16935217697, 
    4755.73309501383, 4560.54645306479, 4281.42897203839, 4002.54091697247, 
    3721.27612304688, 3517.51004318523, 3596.6220612458, 3848.54155667167, 
    4209.41471938769, 4527.88901094197, 4796.56769221631, 5021.14054084063, 
    5199.81641490173, 5323.43922904426, 5394.66730030818, 5382.72491373307, 
    5308.1694774406, 5203.66697922231, 5126.4073229999, 4994.89117254691, 
    4902.4983712602, 4819.10198726848, 4760.91881194588, 4667.27467076735, 
    4502.50539125443, 4256.58131759368, 3975.92038408034, 3757.41747524957, 
    3595.08453826119, 3482.17687430278, 3394.42936943071, 3313.12184463482, 
    3076.1248387077, 2578.1217578457, 2049.34831446174, 1081.54722857398, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 1120, 
    1120, 1120, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 1838.97649596933, 2835.60827823942, 3172.90666787411, 
    3470.49581001404, 3635.25043767152, 3631.97995520467, 3564.78444780552, 
    3463.76519768788, 3361.94043614012, 3306.09500676941, 3202.58497940885, 
    2901.75221911721, 2319.73714776217, 1457.34589636405, 518.736629311704, 
    220, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, 1438.10453256885, 1624.06730079275, 1668.96603338121, 
    1603.41606004546, 1542.80151592839, 1499.13019461423, 1483.25536628064, 
    1371.5613732546, 989.388284282327, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 200, 200, 200, -0, -0, 529.644737532233, 769.392803552175, 
    1142.33014381355, 1673.70716486242, 2210.69268165411, 2594.46067712792, 
    3019.56634683276, 3024.87799954859, 3024.87799954859, 1750, 
    2493.18043927741, 3293.74054183176, 4357.68729126756, 4865.3741469714, 
    5132.25230093171, 5205.43101126826, 5298.49680869563, 5456.85886172462, 
    5500, 5500, 5500, 5500, 5500, 5500, 5149.04343848353, 4894.46810080493, 
    4801.99371904108, 4765.13356703698, 4758.08496382722, 4527.89068240543, 
    4249.56178985823, 3747.04956679511, 3527.03914811408, 3419.3606295086, 
    3387.2978515625, 3844.46884320872, 4472.7961844418, 4757.9867867512, 
    4849.04506135152, 4851.52610453564, 4946.07398654934, 5083.99498581746, 
    5269.82887666949, 5394.45278685228, 5378.83880991895, 5351.75128597706, 
    5271.5545899935, 5207.5738065914, 5178.5908740982, 5047.94360552501, 
    4893.99536029108, 4819.86727614898, 4948.58746082099, 4865.00311145343, 
    4974.93478854665, 4939.60821785119, 4914.58627896758, 5066.16031687674, 
    4963.63561353381, 4623.44261527941, 4118.55991093807, 4021.8546454858, 
    3831.74441800432, 3808.6356057652, 3728.01898233552, 3787.66226256928, 
    3993.80519838615, 4179.68273450409, 4270.09289803483, 4286.2426297535, 
    4453.30390076888, 4553.65407129975, 4544.17843869935, 4419.39777289637, 
    4265.3299316231, 3940.11649356671, 3969.64095854422, 3969.64095854422, 
    4081.49291857824, 4213.35277742997, 4558.94766644972, 4873.60297665893, 
    5115.53620529239, 5237.06641638715, 5255.28186273466, 5238.09290937788, 
    5185.79595627425, 5067.67272395344, 4910.88356251315, 4640.90020911465, 
    4240.78443184887, 3998.57093007234, 3938.53859965485, 3785.16965325578, 
    4527.16129419376, 4901.90755509388, 5133.05376320405, 5266.37071184148, 
    5332.1628747131, 5367.01576884044, 5383.99015082179, 5382.67301265143, 
    5385.31022902594, 5396.93368937005, 5417.8377016733, 5429.15710716779, 
    5436.10782844557, 5445.72568561285, 5418.13630940164, 5361.26461187463, 
    5293.62513549889, 5252.90677177315, 5231.32451205166, 5221.21634110566, 
    5204.38022642608, 5185.03476971507, 5124.31527871197, 5054.94127203752, 
    4978.28977540481, 4891.689773732, 4764.1635758297, 4677.10126740877, 
    4546.67833873783, 4388.38651816804, 4294.18216905883, 4238.59074681248, 
    4163.92461100831, 4105.50418811707, 4043.45059116048, 3971.99957484873, 
    3915.79193481168, 3850.48396639677, 3759.70112106726, 3670.12185603939, 
    3574.98008312386, 3469.58351759463, 3345.8716800008, 3207.86973417009, 
    3178.79671826384, 3225.03356313847, 3230.90243845959, 3123.99238841974, 
    3030.96383105557, 2857.73362143854, 2345.30477155248, -0, -0, -0, -0, -0, 
    -0, -0, -0, 1252.98664018921, 1252.98664018921, 916.045085804303, 
    567.702801697506, 100, -0, -0, -0, 1450, 2025, 3605.48577657099, 
    3708.59949796344, 3495.20937032203, 3496.29436187458, 3337.08116852871, 
    3027.82192117386, 2758.41088867188, 2409.66088288634, 2139.56463702486, 
    1900, 1900, 1492, 50, -0, -0, -0, -0, 3411.11005155238, 4055.67803407735, 
    4342.99704217094, 4342.99704217094, 4121.15725951012, 4282.31880667819, 
    4711.24012772152, 5043.21552264606, 5087.34450649037, 5411.63769009334, 
    5420.34052772997, 5409.14631330518, 5341.79157989875, 5207.51398840714, 
    5101.4450124346, 5015.53432192036, 4903.48809271844, 4787.13365122375, 
    4606.89818572645, 4339.03602268082, 4049.95941678685, 3741.39208726981, 
    3496.86639152958, 3532.31433477508, 3805.48232324858, 4139.74598815752, 
    4512.46779581544, 4793.8139518443, 5017.38353476452, 5204.05284375644, 
    5353.66508835796, 5473.86426802929, 5444.78782148894, 5361.20934212747, 
    5232.13062903418, 5106.07583304466, 4995.56631225873, 4877.51568928711, 
    4803.87550393207, 4761.41220248921, 4704.07114841817, 4619.91514574319, 
    4445.29636481091, 4237.10079538705, 4048.60817787034, 3902.47230445226, 
    3753.1447048037, 3579.99996477992, 3387.44110786267, 3041.58951731484, 
    2506.83537811133, 1888.9850411245, 1081.54722857398, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 960, 1120, 1120, 1120, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    2414.81984229493, 2963.41221211363, 3210.14527338718, 3494.97834217517, 
    3520.33112717251, 3454.30014302387, 3337.57957179841, 3208.27907215275, 
    3116.26409095566, 2918.31688228672, 2548.35330007701, 1838.55198697508, 
    1012.7516976263, 518.736629311704, 220, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, 60, 1142.5, 1101.54602050781, 1061.9, 1008.6, 
    993.3, 90, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 120, 170, 
    170, 50, -0, 80, 100, 180, 1028.5, 1463.4, 1812.1, 2249.1, 2526.9, 
    2537.4, 1900, 2686.1, 3549, 4542.3, 5500, 5500, 5319.6, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5160.8, 4836.8, 4764.2, 4716.7, 4668.9, 
    4426.2, 4102.9, 3621.5, 3522.8, 3452.2, 3615, 4131.8, 4626.6, 4807, 4925, 
    4998.1, 5148.2, 5240.2, 5344.1, 5500, 5500, 5093.1, 5019.8, 5056.3, 
    5056.3, 4881.7, 4813.4, 4779.07568359375, 4857.2, 4989.4, 5112.6, 5500, 
    5159.8, 5247.5, 5176.9, 4957.9, 4579.9, 4355.3, 3981.9, 3765, 3697, 
    3651.8, 3844.6, 4054.4, 4249.9, 4425.5, 4660.7, 4848.5, 4865.7, 4783, 
    4636.3, 4367.2, 4260.7, 4165.5, 4165.4, 4261.6, 4520.1, 4758.7, 4925.3, 
    5018.8, 5033.4, 5003.5, 4910.8, 4788.1, 4621.9, 4368.1, 3969.5, 3560.3, 
    3522.1, -0, 4554.3, 4897.4, 5130.2, 5261.1, 5327.2, 5364.7, 5384.2, 
    5389.5, 5394.8, 5413.4, 5500, 5500, 5500, 5407, 5363.7, 5297.1, 5243.9, 
    5213.7, 5170.4, 5195, 5173.9, 5130.2, 5058.7, 4981.8, 4890, 4826.6, 
    4730.2, 4625.2, 4517, 4403.8, 4304.5, 4237.7, 4170.5, 4115.9, 4054.7, 
    3978.3, 3930.3, 3869.6, 3790.3, 3700.5, 3614.8, 3511.6, 3360.5, 3196.4, 
    3115.9, 3089.9, 3049.5, 2918.4, 2787, 180, -0, -0, -0, -0, -0, -0, -0, 
    -0, 70, 2003.52704338302, 2003.52704338302, 1288.97157337876, 
    1075.02088299144, 100, 40, -0, -0, 1575, 1935.05359591651, 
    3605.48577657099, 3605.48577657099, 3495.20937032203, 3495.20937032203, 
    2992.23551585628, 2367.10580247701, 2072.47117008038, 1741.74447098971, 
    140, 0, 0, 1492, 1492, 943.379565778301, 1196.61395212028, 
    2696.29593328518, 2952.64663076228, 4082.2, 5122.54675447961, 5500, 5500, 
    5500, 5500, 5500, 5271.6, 5293.7, 5452.2, 5401.1, 5345.8, 5314.6, 5238.9, 
    5162.5, 5085.1, 4964.6, 4821.6, 4633.9, 4380.7, 4101.2, 3791.8, 3540.8, 
    3501.5, 3756.2, 4106.6, 4472, 4786.4, 5031.2, 5228.3, 5381.8, 5500, 5500, 
    5403.9, 5260.2, 5107.4, 4987.3, 4870.2, 4821.4, 4829.7, 4856, 4819.7, 
    4700.1, 4538.2, 4373.1, 4217.5, 4042.3, 3834.1, 3567.4, 3112, 2470.8, 
    1668.1, 170, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 960, 960, 960, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 395.982425581927, 2614.3, 3070.6, 3273.1, 3376.9, 
    3311.3, 3178.1, 2983.3, 2764.2, 2513.2, 2095.2, 1118.2, 100, 60, 60, -0, 
    -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, 615.957588262645, 588.490073445489, 
    580.953491210938, 517.996999594479, 503.4209622033, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 50, 50, 50, -0, 80, 100, 180, 
    383.320001348053, 716.033275928036, 1029.69196811173, 1478.68884277344, 
    2028.84029219589, 2050, 1900, 2878.9808965304, 3804.33262430747, 
    4726.93538898381, 5257.40270676689, 5454.20568640249, 5433.73874158606, 
    5346.39143411473, 5356.069399499, 5500, 5500, 5500, 5500, 5500, 
    5487.63695752185, 5172.57376322814, 4779.07571895829, 4726.4824092735, 
    4668.35398567573, 4579.67055776659, 4324.49663005549, 3956.17089331384, 
    3495.99338770107, 3518.63589134862, 3485.0443947249, 3842.79620151924, 
    4419.18185522252, 4780.48294191651, 4856.03812617821, 5000.95390174158, 
    5144.62097498661, 5350.2586422269, 5396.31797260809, 5418.41396986425, 
    5176.63735682973, 5155.30072241337, 4834.39506524005, 4768.08822969502, 
    4795.87949637238, 4934.06795469237, 4715.36379305661, 4732.73123216901, 
    4722.57966926179, 4765.80267180837, 5113.89239765326, 5250.27428069974, 
    5228.44572840981, 5404.9344406022, 5428.79226097062, 5390.26330020859, 
    5292.39651166101, 5041.31443813953, 4688.75146813394, 4132.04400796249, 
    3721.27612304688, 3665.92337521039, 3515.98167277707, 3695.45796098168, 
    3929.17165579643, 4229.67239683302, 4564.660118161, 4868.07942580224, 
    5143.41858983545, 5187.2424974519, 5146.69912043728, 5007.18095939998, 
    4794.35215023397, 4551.68308865095, 4361.27636128503, 4249.35010743988, 
    4309.79051949711, 4481.35181075879, 4643.76557221843, 4735.1180672415, 
    4800.55390639186, 4811.51244377611, 4768.82443246554, 4635.76044531868, 
    4508.60290391542, 4332.89153744089, 4095.2000824118, 3698.27774296668, 
    3121.96360977047, 3105.64634900107, 3919.99034222066, 4581.44328002128, 
    4892.7936157088, 5127.40161870053, 5255.92672988864, 5322.31391504282, 
    5362.38122853939, 5384.43821736791, 5396.35231356534, 5404.38246601009, 
    5429.91452924955, 5464.29089069574, 5467.47436658749, 5417.37048317168, 
    5368.34255733673, 5309.27354040662, 5232.91255588093, 5194.14136622527, 
    5174.42887185671, 5109.50751732772, 5168.75720682689, 5143.41858983545, 
    5075.35341754447, 4993.0343149955, 4908.57553728528, 4801.67340842337, 
    4761.44306418605, 4681.34025903328, 4573.37278606761, 4487.35724069618, 
    4403.8, 4314.87822923518, 4236.82863618165, 4176.99028749994, 
    4126.29456405715, 4065.89147763595, 3984.62943595572, 3944.7390150541, 
    3888.64396798146, 3820.8897521004, 3730.93497250076, 3654.63381634009, 
    3553.6543597008, 3375.19532150199, 3184.83585668101, 3053.09172898444, 
    2954.66819082651, 2868.14576315477, 2712.75358078737, 2543.03849568098, 
    180, -0, -0, -0, -0, -0, -0, -0, -0, 1682.81269153196, 2232.08986350108, 
    2318.75324335053, 1982.80625575353, 1417.97666175447, 766.624765526889, 
    431.797815176131, -0, -0, 1575, 1766, 2758.41088867188, 3141.49507716983, 
    3220.59702967091, 3065.78548661781, 2904.3989830899, 2367.10580247701, 
    2095.33591905228, 1580.9730681579, -0, -0, 1587.81680926245, 
    1912.85780626498, 1912.85780626498, 2593.30125626634, 2588.10940483739, 
    3265.37592741643, 3987.03167792743, 4753.34781405549, 5122.54675447961, 
    5415.53460013457, 5500, 5498.77831658949, 5500, 5500, 5500, 5500, 
    5492.74640301772, 5381.76502652489, 5282.54240676965, 5287.49610086327, 
    5270.2018428692, 5223.48756162596, 5154.57678276071, 5025.77428504109, 
    4855.96665354157, 4660.85285569128, 4422.42076274021, 4152.36215982994, 
    3842.20534426653, 3584.68702156378, 3470.77780538537, 3706.8396772147, 
    4073.46181816253, 4431.54000014394, 4779.07571895829, 5045.10784185514, 
    5252.55404825926, 5409.9383499533, 5500, 5500, 5446.61023459858, 
    5288.306029562, 5108.64324410236, 4979.06240401962, 4862.79346165487, 
    4838.99004535334, 4897.9207067547, 5007.95102538448, 5019.444098968, 
    4954.94380851679, 4839.23507941622, 4697.5790591465, 4532.48973884309, 
    4331.51600455864, 4088.20750858406, 3747.26586721742, 3182.3810921326, 
    2434.8540238458, 1447.17298792799, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 700, 700, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 2265.18296560267, 
    2931.03032835508, 3051.19229219072, 3233.39942891465, 3168.30713527787, 
    3018.61525880215, 2758.41088867188, 2412.11758378817, 2108.02092963711, 
    1642.12574567629, 397.897285337326, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, 220, 243.128140707691, 
    243.128140707691, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 130, 210, 337.38678413084, 569.291861411153, 
    897.941301692752, 1344.65279406825, 1650, 1650, 2831.95305899077, 
    3912.83913846027, 4587.5871318631, 5115.72675009114, 5320.04024773628, 
    5391.0412339335, 5374.25572780683, 5299.26702762467, 5404.45360643337, 
    5485.104423832, 5500, 5490.49769021138, 5418.128147909, 5234.74466767107, 
    5051.21620317841, 4816.90280062366, 4718.06204654026, 4634.43545316812, 
    4434.75639095706, 4100.05650103077, 3662.68170867606, 3502.27996383427, 
    3574.2133861148, 3911.60084290518, 4606.39115667572, 5096.62086450967, 
    5159.27120738877, 5201.81478915991, 5247.43606998025, 5290.04536055634, 
    5362.09143687429, 5354.19183334302, 5326.90976148237, 5186.8260136923, 
    5096.0722872975, 4987.39142593612, 4966.01914867365, 4884.47041730541, 
    4722.3427422077, 4743.26488224897, 4731.67590743849, 4828.45120736322, 
    5026.51363740709, 5306.75023287157, 5479.57443226787, 5500, 5500, 5500, 
    5500, 5500, 5312.17711560217, 5042.75407658872, 4600.74749820307, 
    4128.59247124834, 3893.60395971444, 3968.81636066542, 4026.51440716615, 
    4250.94376144902, 4621.06155004104, 4932.457540361, 5161.87726095317, 
    5342.14904425672, 5371.89044979256, 5330.80200844498, 5177.60575229994, 
    5001.90835600152, 4787.28990069114, 4628.05431500853, 4555.91770472969, 
    4495.10067082505, 4393.42250112511, 4393.42250112511, 4473.96575251901, 
    4494.97601589053, 4482.06168374899, 4479.5824498379, 4387.55136699752, 
    4291.00427036497, 3974.59352956093, 3661.35024422198, 3594.11508060837, 
    3567.81545289294, 3886.35654259379, 4238.95348570643, 4556.10785638462, 
    4888.29441057982, 5155.85386966219, 5260.81710336688, 5344.43196939222, 
    5366.2954958725, 5351.88804430719, 5372.20889399838, 5411.70971981514, 
    5445.46377338794, 5440.75823845869, 5422.78086186214, 5357.89148249729, 
    5307.93160430182, 5240.57979654558, 5172.05228410379, 5129.74043259336, 
    5104.63766859511, 5093.66449145992, 5096.2059966317, 5053.36768939552, 
    4997.92423785204, 4904.26120909517, 4814.3391567194, 4755.5091896856, 
    4690.61628533373, 4596.14192897698, 4494.86194863145, 4403.76222300752, 
    4322.20085359265, 4242.90749327747, 4200.66450931708, 4148.68637070239, 
    4105.99546049646, 4065.89147763595, 4010.50847482137, 3972.53992302803, 
    3911.53780589494, 3858.35177522076, 3769.4559627208, 3687.89276940729, 
    3527.96168859013, 3229.84243547455, 3028.6192429656, 2837.05786008105, 
    2733.67442905946, 2565.7011309992, 2400.53580040285, 1872.69057023415, 
    -0, -0, -0, -0, -0, -0, -0, -0, 1294.90651610182, 2002.05814179379, 
    2526.99224896073, 2637.02709425579, 2637.02709425579, 2016.93197832816, 
    1295.40088498044, 845.497158182377, 479.673847704771, 392.249365634216, 
    1575, 1766, 2039.65292999982, 2224.52709476069, 2209.82712039385, 
    1935.05359591651, 1736.04060688653, 1553.28890800224, -0, -0, 0, 
    899.64290562965, 1567.70525704551, 2041.38286724911, 2368.78820137174, 
    2903.39842204372, 3329.6983367456, 4140.30814486036, 4719.98322905273, 
    5147.78571583169, 5447.79148603634, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5454.36236509268, 5413.86010536901, 5388.92461110865, 
    5351.93463435434, 5268.47130767316, 5132.55969031092, 4948.20283753449, 
    4742.06907111641, 4510.13290104209, 4201.10038303074, 3886.34477764268, 
    3620.57706213077, 3495.23939239972, 3662.52539803985, 4014.47085247991, 
    4388.77659737239, 4723.47261586103, 5007.81583692386, 5232.80804455445, 
    5415.71157239369, 5500, 5500, 5465.1898083533, 5333.7200473915, 
    5227.38790557537, 5127.10364752949, 5054.89441149173, 5072.79149217603, 
    5143.41858983545, 5219.59754179446, 5224.7706441314, 5162.79194009671, 
    5056.31299986824, 4917.31214755645, 4748.27144071311, 4538.62306207064, 
    4271.56841154652, 3887.84055895452, 3275.05437355317, 2527.62442033008, 
    1630.7446304829, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 440, 440, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 2814.21580717198, 2939.94816795681, 
    3030.53881131602, 2953.0914599049, 2744.06343721775, 2409.82714139537, 
    1968.8209235301, 1541.18059616368, 997.956164319738, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 160, 
    294.462890625, 483.353326067035, 663.123067216661, 663.123067216661, -0, 
    2527.2555456303, 3701.00466366145, 4282.5772953884, 4720.62890509443, 
    4916.20956915841, 5119.51454112734, 5225.03738709539, 5180.4396701313, 
    5228.17026741494, 5194.68547444787, 5215.44026104536, 5150.88141900612, 
    5079.13831953717, 4853.46336099916, 4893.42544516645, 4818.95363659772, 
    4722.1096451692, 4592.7309600614, 4263.03224325606, 3853.61287720759, 
    3428.13454370847, 3411.99618904814, 3837.42149899852, 4509.14861378573, 
    5239.51756275973, 5469.1937772164, 5500, 5396.99443064762, 
    5409.27902236899, 5403.58490435225, 5384.80042837547, 5284.21854693643, 
    5143.41858983545, 5164.80441900257, 5105.92512478391, 5120.82085948103, 
    5091.2345614053, 5097.08833762814, 5006.27573743272, 4969.18053117878, 
    4880.08066842642, 4970.92000182487, 5244.48797897039, 5487.57341619208, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5360.92360927813, 
    5038.63949688782, 4766.52068481739, 4470.91112620524, 4579.38975925113, 
    4753.61288382633, 4921.18732836822, 5064.16919983681, 5238.84210710979, 
    5385.57960318962, 5427.95243950157, 5385.90358130139, 5285.73422791572, 
    5161.91857843037, 5004.92568239438, 4824.40173076426, 4695.44315977317, 
    4585.79940418649, 4471.01940194952, 4342.76293489239, 4271.10919654545, 
    4181.19755138833, 4252.48961168686, 4227.54841029466, 4212.53712195527, 
    4109.25843629588, 4107.92556258483, 4127.75313693337, 3986.36491957997, 
    4069.02318845025, 4065.89147763595, 4139.79489735873, 4327.01671339979, 
    4620.59350605132, 4946.15166252547, 5151.01436190436, 5304.3877461846, 
    5362.2873483344, 5366.34259482532, 5367.05849022907, 5376.7136028956, 
    5407.79005436771, 5405.66113339088, 5378.91191081007, 5346.12987108775, 
    5282.81500193214, 5223.04703994679, 5149.49860523745, 5085.98269758974, 
    5051.31651892919, 5004.58543398444, 4995.51200967309, 4989.07725288177, 
    4957.48950148863, 4899.28514475693, 4825.9519383145, 4757.95650892065, 
    4701.79205845043, 4620.78788484811, 4513.48832197358, 4374.91385017379, 
    4312.70324183119, 4218.62875218397, 4184.34860914858, 4172.56187411291, 
    4133.7120977101, 4106.38095583811, 4073.78859253099, 4033.59243985709, 
    3988.55183447122, 3922.84115194424, 3875.42516538882, 3790.32976944914, 
    3639.73709178269, 3388.25576624049, 3076.99138541792, 2689.28024002651, 
    2362.74459947588, 2242.18451503791, 2251.07043846906, 2020.63983158922, 
    1541.71495187922, -0, -0, -0, -0, -0, -0, -0, -0, 1363.00854978339, 
    2118.81533817431, 2680.79249869745, 3122.33778593306, 3140.94292805273, 
    2791.40332945379, 2157.62783253051, 1478.68884277344, 958.204649103509, 
    747.570306540003, 1575, 1766, 1777.96959778234, 1869.08833649555, -0, -0, 
    -0, -0, -0, 382.542757094631, 562.70299923438, 899.64290562965, 
    1603.04486246531, 2243.67548544181, 2915.42217309162, 3758.54177660607, 
    4345.6959150993, 4817.37532568306, 5101.74732796019, 5348.82978242167, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5460.1948490601, 5371.70993748082, 5218.64699103968, 
    5040.03527847818, 4822.60214749124, 4575.55563426316, 4273.86149350807, 
    3954.89326814363, 3676.41075207103, 3519.48037756601, 3638.79619433709, 
    4000.64399197937, 4372.9672379494, 4685.69183746681, 4959.78295744766, 
    5189.59908332579, 5366.93635963706, 5492.3933367049, 5500, 5500, 
    5474.19758337288, 5418.51046875777, 5364.87739597568, 5330.09537187972, 
    5349.75451128321, 5384.10517108612, 5411.67812525665, 5385.45028107325, 
    5307.37170362509, 5188.78180073235, 5051.34329248515, 4875.54377523976, 
    4652.03837831376, 4365.61086671214, 3972.58248492119, 3373.62068139006, 
    2647.00991711195, 1764.17004203156, 1017.00931675316, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 90, 90, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    2698.19068573416, 2839.48086203287, 2817.6282164014, 2645.4649904705, 
    2342.12778557711, 1998.12089995237, 1524.46026246316, 1010.08127328682, 
    650.715690452218, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    253.361404418945, 346.353315645489, 346.353315645489, -0, 0, 
    2838.05986273314, 3241.43072512391, 3563.04857523682, 4016.95019383597, 
    4555.15611342312, 4895.35426495372, 5001.26812444909, 4910.72263796803, 
    4767.71358927335, 4635.41910908366, 4543.29699007952, 4498.29400159493, 
    4647.68921366696, 4753.2691119817, 4700.74361418218, 4754.7458546221, 
    4571.46348337546, 4145.11275256175, 3581.42218783762, 3067.47239076581, 
    3387.2978515625, 4182.49406325869, 4682.64350502973, 5327.09052804218, 
    5500, 5500, 5440.09956204778, 5454.2850089187, 5325.70487303682, 
    5323.72206027581, 5167.83249626458, 5074.06099628222, 5217.56605669813, 
    5289.65663803313, 5326.28583148684, 5149.31249414916, 5207.00593512346, 
    5080.7316374673, 5165.98339180339, 5143.41858983545, 5127.12931167995, 
    5412.18434564344, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5445.99154667536, 5253.92832294059, 5201.30979617825, 5230.38675622809, 
    5292.92952812153, 5379.68343601606, 5432.88140976221, 5480.38356428812, 
    5484.71051347694, 5431.04392878877, 5312.05813498497, 5128.64454953447, 
    4955.93426363363, 4748.98540732335, 4554.41056203977, 4487.28061269262, 
    4332.04027280123, 4208.89830239238, 4107.77235036774, 4041.39143182335, 
    3836.26424760194, 3909.79974301442, 3754.0186501404, 4093.33514804691, 
    4166.96488097987, 4235.42089605154, 4382.0405333897, 4378.32168113366, 
    4331.6351276405, 4319.11791221846, 4367.10795488745, 4530.7425989304, 
    4728.06009263916, 4967.50016156566, 5189.7780636638, 5329.85962579786, 
    5369.84663128668, 5361.88319492535, 5343.30121032628, 5335.32503612685, 
    5329.75545925888, 5318.74388407673, 5277.06290871201, 5216.06445072708, 
    5143.41858983545, 5070.45904698156, 5037.52708169728, 4996.32292357854, 
    4926.07338277115, 4909.65232078179, 4878.56433443683, 4839.46254945775, 
    4851.49755416648, 4814.99803789371, 4757.49214207149, 4696.30503073466, 
    4639.4834823037, 4576.0176020516, 4468.98288371162, 4352.59971416305, 
    4308.91566015912, 4256.55459248428, 4224.81072531513, 4199.35112131078, 
    4158.30918076206, 4119.33038900065, 4084.49486153219, 4049.70161250383, 
    3988.24844343592, 3917.63342240474, 3855.00565555748, 3750.17419383817, 
    3508.18952293575, 3182.85688483383, 2644.9161970204, 1901.47933803023, 0, 
    1613.3515904742, 1613.3515904742, 1493.34795492403, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 1166.34234216907, 1979.39684343851, 2669.92178795707, 
    3232.17939917151, 3261.51385714714, 3261.51385714714, 2933.61012444167, 
    2466.66776221529, 1750.63576409258, 1766, 1766, 1766, 1953.50267444796, 
    1943.5430469766, 1350, 1050, 725, 725, 725, 725, 723.458091322732, 
    1169.381771803, 1891.860826575, 2928.86203462537, 3966.22812861897, 
    4588.32719089546, 4962.2976313046, 5243.08041640052, 5430.50125558659, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5437.36745329945, 5305.42215228244, 5144.17476354817, 
    4913.87086921985, 4643.12110507239, 4328.76882284242, 3994.9240626734, 
    3709.91337222924, 3575.48380666995, 3691.4028177989, 3981.11990026654, 
    4295.5881869399, 4613.74861473268, 4848.78532770921, 5071.37439563568, 
    5255.81225577912, 5420.85524853626, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5464.74936984638, 5363.44497755664, 5244.96529673743, 
    5113.59549083337, 4943.20719313949, 4718.06448095538, 4400.84747301501, 
    3999.41640315845, 3442.53861307656, 2746.82181905041, 1939.40585839743, 
    1154.1565765561, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 550, 1935.05359591651, 2629.68394506281, 
    2700.94699207672, 2661.25234174078, 2448.32131160106, 2179.23838399817, 
    1655.37570446407, 1025.44981546988, 640.130707482274, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 120, 120, 50, -0, 1454.71839500902, 1814.26640540757, 
    1935.05359591651, 2356.95033997088, 3065.78548661781, 4408.9309537187, 
    4408.9309537187, 4396.0340291112, 4348.28311229276, 3911.7656579755, 
    4276.79448339938, 4267.45747236377, 4443.60556552068, 4685.17668708661, 
    4672.76367341456, 4672.76367341456, 4535.43592106507, 4104.06017346922, 
    3326.49188102549, 2840.70704327195, 3275.67806565253, 4182.49406325869, 
    4682.64350502973, 5192.39907638404, 5453.62234873272, 5470.28223753399, 
    5414.87438767584, 5416.21984486357, 5364.37449117547, 5392.80711209425, 
    5185.12344951225, 5327.50597686616, 5253.70648887758, 5500, 5500, 5500, 
    5500, 5445.07718732309, 5399.77093810243, 5260.2100148076, 
    5419.31500436089, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5433.04316034698, 
    5286.49438800183, 5154.00435757885, 4968.77512825792, 4779.07571895829, 
    4480.39522033957, 4277.63479606111, 4240.68851460778, 4096.76319448118, 
    3922.49122516449, 3475.90556876472, 3387.2978515625, 3853.8611271057, 
    4148.77960081076, 4392.31369986562, 4498.59842082107, 4531.33331909932, 
    4527.99127800172, 4538.97401443695, 4566.31232957134, 4606.65542951707, 
    4588.06309114615, 4613.94091886738, 4698.86344947181, 4877.28704639783, 
    5086.09297656207, 5253.72878474439, 5350.68724078472, 5368.99987450881, 
    5363.63733523783, 5339.27557175645, 5301.24692764708, 5252.02072277864, 
    5182.67535004869, 5111.53629039666, 5040.1948658405, 4960.4118196831, 
    4869.8174164645, 4849.90077618417, 4842.38753802309, 4822.56882074634, 
    4790.58002789267, 4745.64756804935, 4698.53772556337, 4727.54682362154, 
    4708.44512416868, 4688.59664638703, 4644.66536766287, 4619.14943386117, 
    4537.9640526432, 4456.60048299223, 4388.82262365625, 4328.58980830466, 
    4299.26474148063, 4243.97435123991, 4233.82435771996, 4177.57399865357, 
    4142.06336437323, 4075.40240865108, 4041.31901875998, 3973.69701162069, 
    3894.45156985319, 3787.38329815986, 3606.57384049254, 3324.21337322215, 
    2888.03433996156, 1810.69215524477, -0, 1084.89265375268, 
    1258.58954725464, 1258.58954725464, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 849.406337366883, 1609.03668898236, 2535.02321027102, 
    3046.31737924758, 3353.76970257869, 3367.83842886924, 2934.2692655717, 
    2992.41248581368, 2711.43833897442, 2321.554024514, 2065.30985669093, 
    2362.54306311021, 2393.2414512705, 2004.8589974874, 1350, 1050, 725, 725, 
    725, 725, 984.384893874752, 1607.82027315826, 2594.14006092537, 
    3861.49067175658, 4646.2098511191, 5094.05396128603, 5361.55184393308, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5466.96875717598, 5357.25636868183, 
    5146.80188254949, 4931.8935363094, 4702.83431887345, 4367.43087740036, 
    4002.28238333452, 3658.0376399383, 3536.29234831545, 3677.67339380982, 
    3877.59444043501, 4186.5217297236, 4462.42788905638, 4706.27652390386, 
    4909.82517234916, 5110.7396448748, 5290.33616398043, 5428.56030560264, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5441.97248033712, 
    5361.18544682757, 5246.52278298365, 5132.39306222547, 4977.88895173951, 
    4761.42232545537, 4449.82128318751, 4044.14785200989, 3522.63891345099, 
    2886.91707803041, 2313.84190817368, 1466.64222434371, 946.697003662581, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, -0, -0, -0, 
    543.685815962427, 543.685815962427, 1935.05359591651, 2099.11988533156, 
    2078.12587358242, 2144.19445271096, 2037.14581171507, 1909.15491922942, 
    1494.17101832261, 705.375280893213, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 50, 90, 170, 708.028137663733, 1101.54602050781, 
    1478.68884277344, 1628.42738007182, 1716.61708354511, 2690.6068224277, 
    4065.89147763595, 4334.80885140077, 4092.57435273921, 3890.24368219647, 
    3768.06146287676, 3863.22450696005, 4250.72107120215, 4250.72107120215, 
    4765.88167919095, 4706.63340322074, 4600.36146813833, 4001.23123349367, 
    3124.25908818257, 2940.43947333479, 3065.78548661781, 3634.11519420264, 
    4373.32867966005, 5094.68127969617, 5094.68127969617, 4996.10970298439, 
    5184.4655763792, 5500, 5500, 5500, 5480.55706134194, 5366.94478519537, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5433.48334136386, 5292.56704445747, 5107.30464346783, 
    5013.7551650431, 4859.87542221339, 4440.31456315733, 4141.60718152867, 
    3707.90617405782, 3687.27626826911, 3032.98897132766, 3187.25297801123, 
    3104.32321509862, 3534.88946302815, 4278.9971761775, 4403.51916943482, 
    4559.489094461, 4685.86046830051, 4727.17368377389, 4700.38689071824, 
    4648.1225106441, 4710.16495341393, 4779.07571895829, 4805.73751262126, 
    4872.48606343551, 4969.97932752489, 5110.42043183346, 5248.95657210893, 
    5350.82896020045, 5393.23702682599, 5390.85471975478, 5347.72916859008, 
    5292.12782454226, 5253.59345156474, 5165.96098559502, 5103.79635465292, 
    5017.19101665827, 4919.04222658578, 4846.08657826534, 4765.34059159893, 
    4762.26129998763, 4762.26129998763, 4735.85079016666, 4734.90078624572, 
    4700.43430455542, 4685.37882807896, 4657.66058122337, 4628.38027278946, 
    4494.23077591401, 4618.53090025146, 4602.36139609532, 4541.51470135921, 
    4438.06492459607, 4382.86983473999, 4403.57248540015, 4394.21162043642, 
    4290.50809748303, 4244.16048372244, 4163.06840945392, 4114.87079211772, 
    4054.04181015253, 3884.57361783918, 3895.97699235018, 3875.75174900093, 
    3738.90249942298, 3492.68395295446, 3078.9385323114, 2126.33682669641, 
    1101.59687702663, -0, 1063.80305233146, 1017.54041577472, 985, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 495.553629324057, 950.990525108759, 
    1853.60996436837, 2644.86488949539, 2891.78987884444, 2934.2692655717, 
    2962.49563891149, 2931.29124621629, 2711.43833897442, 2532.46529351453, 
    2688.16259252811, 2723.79241932252, 2493.46757975451, 1766, 1050, 1050, 
    725, 725, 725, 725, 1045.7060178942, 2288.9680100775, 3768.28077916148, 
    4381.39460977881, 4966.9555845964, 5291.28554886568, 5434.63454115527, 
    5498.46342714342, 5500, 5484.25862629629, 5437.99647702269, 
    5431.9411302532, 5425.68027447582, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5472.699330535, 5338.63525490882, 
    5155.96445885222, 4936.34413432883, 4695.87005211044, 4428.22289157311, 
    4106.8436290405, 3799.19787249147, 3507.27397402021, 3575.76732696217, 
    3768.87920627536, 3978.22686642523, 4262.95200827403, 4511.23730923776, 
    4731.9010610034, 4969.52264199609, 5127.60480516181, 5287.87167667909, 
    5421.4556783612, 5500, 5500, 5500, 5500, 5500, 5495.96782361793, 
    5411.81963766389, 5337.51955234786, 5221.0985577023, 5201.96039698425, 
    5132.39306222547, 5010.63397583113, 4821.81554245587, 4544.18646984597, 
    4181.77930223827, 3554.5096735072, 3193.09711400127, 2830.77749578042, 
    2153.87076477805, 1119.75151628386, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 0, 40, 40, 40, 40, -0, 543.685815962427, 543.685815962427, 550, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 50, 90, 170, 240.561416625977, 309.700115949049, 
    433.214550151211, 1037.21746170963, 1184.90401825481, 1184.90401825481, 
    2069.15673603546, 3977.51504865436, 3721.27612304688, 4148.30459798986, 
    4641.93218948168, 4627.28038764959, 4581.02722050418, 4138.5666110755, 
    4706.63340322074, 4706.63340322074, 4596.63802945649, 3947.2828866379, 
    3200.70963089873, 2940.43947333479, 2741.65215227743, 4234.79623816193, 
    4234.79623816193, 4864.36688531722, 5273.84370579979, 5478.02837088514, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5460.75948415067, 5416.37768416819, 
    5239.20876918856, 5108.59662581777, 4892.75951864191, 4561.17106936914, 
    4561.17106936914, 4307.78854209189, 4385.6473963492, 4385.6473963492, 
    4373.96977209787, 4332.38181302157, 4195.66411979679, 4065.89147763595, 
    4200.95345430134, 4339.27744788623, 4557.74923313882, 4790.17421855892, 
    4880.10599221706, 4941.58654902576, 4745.79942610636, 4612.08931412022, 
    4692.1933650918, 4870.92120623191, 5097.80356993734, 5143.41858983545, 
    5299.54393487255, 5376.83255203848, 5389.83214466925, 5386.9609100072, 
    5437.15623430912, 5374.66309006802, 5390.32416176826, 5335.28606310667, 
    5235.49819936235, 5143.41858983545, 5060.94183794691, 4953.78887898184, 
    4860.20278673765, 4779.07571895829, 4779.07571895829, 4746.95450986098, 
    4715.05717276483, 4731.56395956589, 4692.51951276439, 4632.74816193669, 
    4576.27024111388, 4541.42804642691, 4552.18805381583, 4511.20386551103, 
    4568.27165251778, 4591.8428158894, 4543.67442822181, 4499.0114652462, 
    4457.58879399485, 4422.49231960914, 4383.7826771438, 4257.80051418926, 
    4224.00627586184, 4065.89147763595, 3961.27758532308, 4028.70077653182, 
    3966.26387465698, 3968.10221385396, 3805.09773243117, 3580.345822392, 
    3355.15054275508, 2817.25440383604, 903.202372644174, -0, 200, 
    358.842227607406, 358.842227607406, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 513.396786309341, 1378.86625986848, 1706.37581171375, 
    1783.96082118797, 1941.91155541721, 2525, 2525, 2617.47380214645, 
    2532.46529351453, 2688.16259252811, 2694.42088391493, 2493.59680075172, 
    786.194940018987, 356.604517382195, 130, -0, -0, 725, 725, 
    1045.7060178942, 3558.81249184459, 4226.83864283473, 4527.02835363683, 
    4934.73968249927, 5166.75284031008, 5365.58217848903, 5468.46711209483, 
    5425.73997822349, 5365.80376369909, 5318.61467748255, 5184.32727517156, 
    5300.79227686046, 5374.06042449425, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5442.65808320394, 5343.37886869309, 
    5215.02829147861, 5001.16121480734, 4785.26818818361, 4554.62450040195, 
    4252.26313535976, 3882.01491896553, 3595.67083316384, 3370.12177491397, 
    3581.80040882705, 3828.58687372342, 4065.97252563399, 4360.59267932207, 
    4621.96482260372, 4843.33191781862, 4978.29345010084, 4990.46556513478, 
    5152.09480386892, 5368.69432659133, 5413.08088233083, 5500, 5500, 
    5444.87372548329, 5346.99512374499, 5266.95913931738, 5158.44330946732, 
    5143.41858983545, 5150.83524074558, 5126.39819761535, 5029.60096887841, 
    4883.84501439558, 4669.87323600178, 4332.09578639188, 3920.05694273283, 
    3542.93338387968, 3276.68673418767, 2989.07003855752, 2281.01743649707, 
    1052.6021094987, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 
    0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 40, 40, 40, 40, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 80, 130, 130, 210, 258.619819757225, 1091.45759632561, 
    1091.45759632561, 761.186687149552, 2168.53254680227, 3721.27612304688, 
    4148.30459798986, 4498.79480658332, 4671.63422504055, 4442.19020711976, 
    4614.25643351469, 4651.93723626906, 4651.93723626906, 4502.45435087847, 
    3313.21924373371, 2867.74369731689, 2867.74369731689, 2395.75572735758, 
    4987.55844482179, 4987.55844482179, 5086.25709241021, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5369.26244336745, 5319.93197884262, 
    5293.39360278955, 5174.13869473714, 4704.75757195797, 4702.76173058714, 
    4702.36779545275, 4377.10252661145, 5131.70947389774, 4997.1725949021, 
    4863.09323791374, 4764.16675529655, 4493.82810334713, 4435.30343589932, 
    4406.84883740431, 4485.0552508499, 4638.21888795583, 4797.40753479764, 
    4980.67585162099, 5006.16268921179, 5029.85841018616, 4221.99630830363, 
    4762.56432235319, 5009.67051417345, 5150.09446168595, 5434.42707381433, 
    5458.48496684221, 5500, 5500, 5500, 5466.27226717777, 5458.26768365846, 
    5348.98783705145, 5363.93213116636, 5254.48763452543, 5121.17018980454, 
    5093.27094962294, 4977.6464436379, 4854.43953988187, 4879.93397503383, 
    4869.85203783955, 4812.87518570671, 4845.00582020524, 4735.60964879411, 
    4735.60964879411, 4712.39546873983, 4627.60915241338, 4568.72025674217, 
    4419.18185522252, 4465.41351635415, 4451.46445272772, 4357.98529411924, 
    4461.1620604958, 4498.22733307034, 4471.94267248149, 4503.43898412141, 
    4425.39504250863, 4390.83572188673, 4287.19301866338, 4265.72860124677, 
    4233.63495227896, 4038.82489724606, 3986.65427142924, 3853.26055307463, 
    3796.02787603325, 3660.5916009633, 3521.32515238926, 3093.22250613401, 
    50, -0, -0, 200, 200, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    170, 735.083559578118, 735.083559578118, 690.06230864761, 
    907.937042598612, 1101.54602050781, 1223.74321593965, 1673.63556022877, 
    2075.34014132633, 2570.78436860381, 2683.96271726195, 1723.56624059178, 
    352.631598590579, 140, 0, -0, -0, 725, 725, 1134.50781640627, 
    3458.98079440547, 4547.02934421378, 4610.43159623756, 4779.07571895829, 
    4992.80991157666, 5336.52659831274, 5471.16532678084, 5437.13518501011, 
    5305.41946926374, 5104.66038595275, 5105.25228847183, 5271.28069253387, 
    5237.05798986722, 5460.36156260551, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5462.23757332069, 5411.42944085553, 5253.13353081636, 
    4942.47609321592, 4781.52711271885, 4472.54120392484, 4290.67005999108, 
    3954.40790753497, 3708.64589582527, 3102.12362495289, 3195.54561423941, 
    3732.39651611362, 4014.84282943856, 4108.40196727582, 4506.01698541743, 
    4657.7181022409, 4779.07571895829, 4925.23550857279, 4987.13681072286, 
    5094.03210275424, 5189.41734380107, 5254.2498349099, 5164.25569893891, 
    5095.8401473569, 5121.37198600958, 5121.37198600958, 5126.52601722084, 
    5126.52601722084, 5228.55190745549, 5172.78123443397, 5048.66913887088, 
    4916.07403923545, 4779.07571895829, 4541.23941136016, 4217.60109401583, 
    3756.68239931936, 3276.68673418767, 2989.07003855752, 2204.8498767428, 
    2225.68862910104, 582.717608576429, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 
    0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 80, 80, 90, 130, 130, 761.186687149552, 
    761.186687149552, 425.785466617812, 2191.85384798669, 3451.50719380881, 
    3451.50719380881, 3902.208732265, 3902.208732265, 4554.67148512565, 
    4554.67148512565, 4439.99924900832, 3801.2956259648, 3284.25886035248, 
    2466.66776221529, 3187.50203223402, 3187.50203223402, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5470.45570974767, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5449.40978225851, 
    5180.58670489665, 5116.07221732528, 5273.80624717664, 5254.76093866463, 
    4759.66290976541, 2666.85344961206, 3700.09372782084, 3450.79160480747, 
    4678.42189698653, 5294.58801717961, 5178.71068978265, 4961.96717246568, 
    4779.07571895829, 4804.50558257091, 4704.40565240338, 4787.82983296497, 
    4874.54429387878, 4981.16716527548, 5074.0436565601, 5074.0436565601, 
    5006.16268921179, 5103.12344031651, 4987.24443976158, 5287.80430132643, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5490.81564207919, 
    5435.63890688355, 5429.17626904116, 5338.36994805244, 5248.954052171, 
    5021.35857233725, 4852.38484874584, 4888.88365661156, 4925.41937427591, 
    4925.41937427591, 4896.68165624002, 4897.78119116183, 4800.47220999118, 
    4811.05235130186, 4735.60964879411, 4608.20061408245, 4581.91441512575, 
    4256.77221410031, 4173.63742047545, 4259.28834051662, 3975.45119585192, 
    4274.56230393198, 4562.86608287282, 4476.18310894635, 4438.60341717844, 
    4473.7878551556, 4446.25127928098, 4352.63059624182, 4288.47788968519, 
    4320.79334883571, 4225.26893329161, 4038.82489724606, 4031.05219900329, 
    3856.27980212675, 3703.30040508766, 3587.72162480898, 3699.4281977897, 
    543.460995719773, 50, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 40, 40, 60, 70, 80, 80, 90, 495.553629324057, 
    1560.57440305653, 1560.57440305653, 640.054220822384, 259.969334952472, 
    90, 40, -0, -0, 40, 757.21070163853, 836.232719608352, 1134.50781640627, 
    4292.5285962713, 4592.43163489512, 4728.55683568012, 4654.28189419278, 
    4802.13116646362, 5290.588482308, 5423.49237798131, 5497.26849604017, 
    5275.03753893143, 5086.04991921922, 5105.25228847183, 5105.25228847183, 
    5079.3403492301, 5239.55877142088, 5456.94686795654, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5459.69704719626, 5397.36393958745, 
    5328.10559776886, 5072.1410423029, 4842.10073299794, 4726.49951891595, 
    4389.19816633122, 4015.18786875292, 3700.56682806799, 3276.55148499328, 
    2973.08820173744, 3421.45661051468, 3752.54555124262, 3844.51072469899, 
    4065.89147763595, 4455.61676134826, 4519.74087547082, 4618.26780950846, 
    4767.9997669222, 4833.72938821926, 4898.60218545016, 4893.21759457718, 
    4726.70120370076, 4823.37898706989, 4817.25159730609, 4879.33395450505, 
    5097.58709447162, 5187.87956525022, 5295.57958100995, 5229.09769426358, 
    5077.14512470421, 4946.77532446575, 4835.93392821747, 4664.89761499337, 
    4384.28742160037, 3964.37741118265, 2278.90947677801, 985.310435888532, 
    2390.40414300927, 2390.40414300927, 1234.35694084501, 180, 80, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 40, 60, 60, 80, 120, 457.436638995133, 
    457.436638995133, 381.207025900257, 968.280578226035, 3451.50719380881, 
    3451.50719380881, 2921.99712859953, 4326.44425777797, 4547.91603828708, 
    4493.5351350664, 4271.69744938501, 3506.61258753717, 2679.21201976696, 
    2481.14037813022, 3704.12954730825, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 3810.09540801161, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 4268.51809268999, 4946.21949950423, 5189.45875378886, 
    5194.35264952418, 5116.07221732528, 5116.07221732528, 4586.87690100807, 
    5234.62900334248, 5408.3225510656, 5439.90815293528, 5366.54498400489, 
    5269.75449997378, 5296.47994038452, 5257.20195182626, 5002.20986462044, 
    4964.7607994457, 5101.24803606542, 5143.41858983545, 5221.86215082407, 
    5204.32073856864, 5270.21906675407, 5352.53929092334, 5357.29519909301, 
    4626.66150618007, 5500, 5442.10695335002, 5481.21686759631, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5356.31707726467, 5373.79773362072, 
    5254.17048484693, 4815.97471991651, 4700.0381198552, 4907.71330962704, 
    4823.52474866296, 4978.86222545965, 5070.05951135519, 5000.51724887375, 
    4956.9453010046, 4930.87482539234, 4779.07571895829, 4642.67247757111, 
    4233.6680213955, 4245.5997145428, 4245.5997145428, 4065.89147763595, 
    4403.5786216881, 4386.06190501498, 4481.06099553392, 4677.70147252486, 
    4608.21661745763, 4511.98262819734, 4426.98218149044, 4257.8420520743, 
    4387.42862497139, 4309.72757977987, 4260.29559987769, 4193.87070523279, 
    4001.19273819045, 3896.38129712542, 3464.770369882, 3216.39132227544, 
    3146.23664453202, 1668.82076305403, 110, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, -0, -0, 0, 50, 
    230, 230, 40, 40, 40, -0, -0, 40, 769.346451300268, 836.232719608352, 
    920.155490936288, 4368.80047847232, 4592.43163489512, 4592.43163489512, 
    4231.17784076216, 5010.34677833567, 5433.68843475497, 5454.36576127352, 
    5330.18868989744, 5242.36593588736, 5165.32351268771, 5086.04991921922, 
    5005.54407801367, 4941.11557825738, 4982.61913451037, 5047.38351221901, 
    5213.06067351008, 5471.03747919457, 5500, 5500, 5500, 5500, 5500, 
    5443.75796481753, 5403.28216615098, 5398.49858988671, 5201.38446675581, 
    5031.75826681908, 4990.74000788849, 4688.85490445163, 4338.30998605763, 
    3988.84734677484, 3690.80419569813, 3666.0494610969, 2992.08811326625, 
    2689.37295790004, 3280.40316942784, 3500.9552948781, 3847.29470732024, 
    3888.30106161791, 4065.89147763595, 4389.00853516062, 4664.11109018134, 
    4675.52357847591, 4563.44193513419, 4642.3920110745, 4616.53202253023, 
    4592.62328997775, 4419.18185522252, 2985.84476066458, 4973.64573723084, 
    5146.75499593097, 5315.39203786521, 5335.09605890279, 5177.58664636368, 
    5042.21440654942, 4882.78283746108, 4744.171118317, 4570.98521933854, 
    4378.10827556442, 4119.94360013601, 3751.58657695638, 3641.53938702883, 
    3009.54983235387, 1402.15791370575, 1488.65332719015, 1488.65332719015, 
    337.896148266657, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 0, 40, 40, 50, 50, 90, 150, 495.553629324057, 
    495.553629324057, 90, 1679.52972118451, 2921.99712859953, 
    4515.77437914091, 4544.11329260969, 4326.44425777797, 3997.32758927277, 
    3997.32758927277, 3178.39513003479, 1759.80757568256, 1570.1704734156, 
    3521.34267244508, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5162.64271951156, 5209.42850650674, 
    5337.72997689525, 5345.82811751425, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5152.41012939708, 4999.56933124315, 
    5054.09855975076, 5089.42691724419, 5076.03942126087, 5076.03942126087, 
    4621.96895337652, 4803.44454604602, 4935.80620900274, 5320.55674269753, 
    5192.90817611579, 5242.58280204114, 5258.3132860105, 5211.39893711188, 
    4531.34798047161, 5383.35914039558, 5312.09875540169, 5438.27108093355, 
    5449.29774851873, 5492.21538584738, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5352.89491639186, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5494.87929720747, 5269.78940217349, 5209.7469464129, 5299.76987257933, 
    5411.9158441857, 5365.87840336452, 5496.29616592046, 5339.96043052678, 
    4982.67609029232, 4997.02540127852, 5083.86447742673, 4728.05403243837, 
    4730.72815881575, 4730.72815881575, 4603.11147968976, 4357.21926708419, 
    4180.39756835179, 4372.91722198772, 4549.87150245163, 4672.00350387515, 
    4425.2509405837, 4710.64930681819, 4575.83895191083, 4575.33092685022, 
    4499.83034192987, 4488.93441861115, 4305.77303087188, 4287.87506271993, 
    4123.79246867012, 4200.2125480588, 4030.42921696512, 3906.2238112085, 
    3966.36551175895, 3891.06849711065, 3646.2931709095, 3010.49334173683, 
    2222.58400988417, 1567.18678192427, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 0, 40, 748.158466361998, 826.63092370477, 
    920.155490936288, 3512.63949136822, 4048.70715668146, 3848.45426115657, 
    4916.98230639748, 5343.92718686525, 5414.97395745251, 5415.44147795045, 
    5319.93440131734, 5206.10797593873, 5143.41858983545, 4989.04205990515, 
    4853.18687837358, 4672.01020068447, 4856.43116858309, 4882.58616228136, 
    5035.68874408436, 5376.33943979005, 5476.71653787622, 5387.97286768633, 
    5500, 5500, 5500, 5458.3287076987, 5500, 5364.14519868137, 
    5395.14427643736, 5097.19948850821, 5071.61284570711, 4822.23751505788, 
    4419.18185522252, 4130.05047199556, 4043.49279222019, 3894.44750721247, 
    3443.53075815251, 2980.75744096045, 2588.06291459658, 3294.15155892356, 
    3421.41438093875, 3614.30313803241, 3650.34889373461, 3864.78044566008, 
    4419.18185522252, 4419.56547970075, 4523.34025506215, 4649.87049496869, 
    4518.39704688123, 4556.83984550192, 4302.82469340023, 2985.84476066458, 
    4675.1352471986, 4939.23677375357, 5335.45571268366, 5411.3731998043, 
    5326.63589161238, 5124.97040770217, 4934.85643017528, 4853.01453984159, 
    4757.20095811883, 4596.37736989291, 4432.18189249813, 4065.89147763595, 
    3621.63866003539, 3009.54983235387, 2138.27858998356, 2120.70711350921, 
    2120.70711350921, 1168.58181957785, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 0, 40, 40, 50, 50, 80, 150, 495.553629324057, 
    495.553629324057, -0, 140, 2347.64323449113, 4658.70917247266, 
    4430.38276135287, 4043.3666157034, 4043.3666157034, 4037.0292233418, 
    3065.78548661781, 1147.43888841087, 1962.02646091024, 4478.01349718842, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5467.25859622689, 
    5500, 5500, 5500, 4848.13995659466, 4193.80411989706, 3962.02788176693, 
    3610.43972832895, 4320.817205232, 5401.80921905009, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 4999.56933124315, 
    4999.56933124315, 4946.94680839765, 5298.01806041953, 5364.13225659414, 
    5312.54850012697, 5151.14742718001, 5248.2638977767, 4935.80620900274, 
    5178.94330366748, 5287.89547347067, 5419.59180818559, 5373.72915342201, 
    4713.86184317215, 5391.7765530756, 5487.41335729049, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5448.00097862827, 5480.78571725452, 
    5060.50697903376, 5493.38088228668, 5460.45406675316, 5500, 5500, 5500, 
    5500, 5500, 5500, 5439.18542180991, 5349.60775117215, 5156.0181903065, 
    5357.92723128805, 5442.12518243701, 5500, 5388.25731834803, 
    5461.73391978873, 5485.50893536456, 5500, 5500, 5181.70152588629, 
    4976.19756801729, 4688.74629983704, 4638.08273602956, 4688.51199101774, 
    4727.20124337939, 4552.84491455234, 4732.03422774582, 4633.77534111483, 
    4606.87928172722, 4602.51440492256, 4526.05397686693, 4506.40475097284, 
    4395.31380092304, 4219.02942414092, 4185.52152047021, 4204.04441856964, 
    4224.09889946603, 4118.34101694137, 4096.1159118154, 3976.37715951696, 
    3938.95203072869, 3915.08391642012, 3409.96777948763, 1649.37443571778, 
    1517.40493584456, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 40, 335.522604658122, 725, 899.074372840564, 
    2715.25457598191, 3092.30794343839, 4368.34332012582, 5114.56477052343, 
    5412.67088493108, 5443.30452610909, 5436.52209222747, 5360.06456812806, 
    5219.48317888596, 5087.80308040875, 4908.91491409218, 4684.96551946354, 
    4420.36154512503, 4548.17335819077, 4711.90028773422, 4784.39790463933, 
    5227.76388566458, 5226.07947700931, 5417.62667054708, 5500, 
    5469.45654447716, 5500, 5500, 5490.52208586754, 5432.20160869515, 
    5468.02550137871, 5097.19948850821, 4965.34031316527, 4830.06480868348, 
    4813.47138576479, 4721.5460595729, 4189.11552903613, 3806.02307925765, 
    3480.98894969224, 3331.94755963062, 2662.26669987456, 2648.84278997312, 
    3297.73918029072, 3419.66282965061, 3403.64810990363, 3772.50342719021, 
    3812.90723834022, 4180.80165736273, 4232.38424616397, 4193.65322524482, 
    4398.18757713531, 4131.9505161422, 4113.27284014808, 2033.18460502804, 
    3993.72621048776, 4939.23677375357, 5376.02217683495, 5438.22406257953, 
    5390.14751726762, 5203.31108129562, 4982.86705962595, 4837.30924925493, 
    4626.43461708798, 4681.80073918165, 4524.43446924658, 4065.89147763595, 
    4393.36978322367, 4129.6327406945, 3138.87149437924, 3342.01660755375, 
    2503.44334290523, 1168.58181957785, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 160, 
    445.999352660532, 445.999352660532, 370.848607337333, -0, -0, -0, -0, -0, 
    40, 130, 1327.38179119433, 1327.38179119433, 812.469668752819, 0, 0, 40, 
    40, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 40, 40, 50, 60, 60, 80, 150, 150, 150, -0, -0, 
    952.454139203525, 977.252984454408, 2841.1344229216, 4043.3666157034, 
    4043.3666157034, 4037.0292233418, 2977.20093318978, 905.427415331652, 
    2027.03687450736, 4588.67186019055, 5500, 5500, 5500, 5500, 5500, 5500, 
    5070.96020963902, 5500, 5500, 5500, 5500, 5365.17637331415, 
    4811.67350364737, 4510.45434029078, 4581.67521103752, 3138.93238018998, 
    2559.12237988314, 3958.57447615096, 5224.3033737235, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5491.65346485113, 5307.88509075293, 
    5321.50007391959, 3291.49582151633, 4946.94680839765, 4946.94680839765, 
    5300.53346945001, 5290.64039341892, 5320.40796833544, 5143.41858983545, 
    5231.79968663382, 4935.80620900274, 5277.1069714994, 5274.47567332242, 
    5327.45398964826, 5009.12431537374, 4791.12619733219, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5351.11212640774, 5061.4366196557, 
    4856.17617982649, 5130.02021021091, 5320.20923918272, 5500, 
    5451.68342984431, 5500, 5500, 5500, 5500, 5500, 5424.73951726343, 
    5429.33034073007, 5418.3405571902, 5355.00357726649, 5490.154419791, 
    5500, 5500, 5500, 5303.32871898712, 5500, 5384.62721031194, 
    5255.97179080715, 5093.42503292241, 5082.91045144029, 5009.03835800477, 
    5037.88708343826, 4853.99515533048, 4788.34123350214, 4542.55552664981, 
    4419.18185522252, 4524.36500391123, 4505.39337371137, 4474.72983085679, 
    4288.61915756879, 4270.04822089267, 4270.04822089267, 3895.5919677285, 
    4298.60646016525, 4334.23506769948, 4334.23506769948, 4204.26490588131, 
    4160.17929924221, 3774.73741611514, 3707.69068154064, 970.336041769536, 
    970.336041769536, 928.924241949538, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 40, 350, 625, 1626.58827909485, 
    3257.191237058, 4368.34332012582, 5114.56477052343, 5337.09705562664, 
    5398.82960692527, 5410.76174841736, 5351.52000242709, 5193.71076202838, 
    5101.76715238234, 4906.25507832382, 4736.95127100806, 2328.44055700253, 
    4500.6419754464, 4683.36710266548, 4583.01592216831, 4653.34982337321, 
    5160.53849096404, 5166.00611698091, 5319.75406755581, 5500, 5500, 5500, 
    5500, 5433.95539977494, 5438.52056938892, 4317.71664000694, 
    5050.86182321678, 4996.22009384942, 4989.97353957946, 4629.08103968976, 
    4172.15970865809, 3975.11060602199, 3814.94330058187, 3451.81298226909, 
    3423.39292631393, 2692.95500097693, 2603.30719410179, 3079.31352513963, 
    3237.96565346693, 3475.59061001256, 3456.33505119562, 3695.19754497184, 
    3828.11586242859, 3924.67809179961, 3694.88917693318, 3594.12508570708, 
    3588.56693904547, 2682.19299911266, 2540.88730261653, 4870.39150213169, 
    5096.93381780119, 5376.41316705556, 5407.55333968837, 5266.72599257907, 
    5132.81544331448, 4831.47431804297, 4045.709830382, 4045.709830382, 
    3584.62744992475, 2223.97957773313, 4317.92449442563, 4374.55151644433, 
    3815.19596108826, 3792.45110812078, 3398.85751626303, 3497.1011209904, 
    180, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 0, 359.039109051824, 1208.10912140781, 
    1794.4470397205, 1840.87507319538, 1035.26562252102, -0, -0, -0, 
    375.368414847542, 1740.25407539853, 2384.42589520022, 2530.12487545024, 
    2650, 2650, 2213.91437577074, 1595.08539089752, 1266.95791675348, 
    1155.36229246683, 1155.36229246683, 908.805143757966, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 0, 40, 40, 70, 70, 60, 70, 150, 150, 150, 150, -0, -0, -0, 
    472.698397477378, 428.807038515461, 2053.13441399311, 2796.69405919677, 
    2796.69405919677, 905.427415331652, 1137.0147741529, 5500, 5500, 
    5431.77802592941, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5391.92884818025, 4437.137198342, 3319.57160336008, 
    3522.35049857784, 4450.56913853549, 5483.61005227974, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 3414.86881756021, 3311.58459987263, 
    3736.16308583393, 3736.16308583393, 3024.50645111369, 2895.00652193514, 
    2895.00652193514, 2813.36953801248, 2500.38416677981, 4704.52177023344, 
    5074.55804153583, 5006.66111122375, 4335.09705172939, 4999.27718787381, 
    5414.91126273124, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5166.87869274777, 5500, 5364.72879982916, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5483.80294700691, 5447.02996019211, 5326.29786161346, 
    5333.66330965034, 5238.92227013074, 5095.1824407412, 5095.62663154154, 
    4998.34663652118, 5009.74090147413, 5039.00175471818, 4730.27531724015, 
    4938.4083646521, 4960.28515948611, 4998.13957041328, 4958.78649491966, 
    4911.32773234208, 4637.96905133617, 4596.47888426957, 4439.74218431627, 
    4378.28326039716, 4408.53490092735, 4379.38991856722, 4240.36384324183, 
    4146.04067521146, 3625.12274099329, 1306.45741483789, 962.84893935623, 
    617.501089981583, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 40, 40, 464.145383636434, 3257.191237058, 
    4226.16060514707, 4688.83664618985, 5117.5516577604, 5342.74717848095, 
    5358.05970704077, 5387.3991500379, 5290.72679534501, 5117.18981914939, 
    5077.80517628447, 4866.94256024976, 4696.50197817043, 4762.31043908007, 
    3869.84372610951, 4315.81630725289, 4541.32464079141, 4671.94828967152, 
    4671.94828967152, 4779.07571895829, 5460.97014686528, 5500, 
    5459.06440010919, 5500, 5500, 5182.39403778142, 4317.71664000694, 
    4996.22009384942, 4996.22009384942, 5126.12063986036, 4677.09608793395, 
    4556.71429717129, 4012.99836049428, 3858.28318974582, 3689.90922045715, 
    3689.90922045715, 3242.17157721654, 2421.25832110625, 2596.63100807026, 
    2724.83768302018, 3173.49036899828, 3271.51929880419, 3310.62806264413, 
    3310.62806264413, 3434.06868469564, 3440.76479761877, 3290.4387064614, 
    2682.19299911266, 2874.01903861248, 4002.24540602273, 4425.11483770539, 
    4880.91629572279, 5201.12044154342, 5383.39270743014, 5342.07501251266, 
    5319.51442523954, 5173.37978600885, 4535.76712949885, 4107.25611177991, 
    3863.92576957812, 3467.57508227944, 3905.77500508155, 3815.19596108826, 
    4194.39150875792, 4309.82843176136, 4344.83908641434, 4367.69650083369, 
    3008.62135438261, 140, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 40, 90, 230, 302.029492921295, 
    359.039109051824, 1650.16416642798, 2276.73607210723, 2617.64440214332, 
    2703.59399301473, 2703.59399301473, 2338.39100696543, 2050, 2050, 2050, 
    2384.42589520022, 2530.12487545024, 2650, 2650, 2650, 2650, 
    2246.96905258671, 1495.41326123443, 1155.36229246683, 908.805143757966, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 40, 40, 70, 80, 80, 60, -0, 150, 150, 150, 150, -0, -0, -0, 
    -0, -0, -0, 398.129436476749, 686.841575071371, 686.841575071371, 
    1137.0147741529, 5500, 5500, 5480.84314236749, 5448.72889284061, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5399.20255493904, 4583.96945020067, 4391.2578033778, 3665.02278694042, 
    3923.01190813782, 4808.14815026151, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5398.9989531454, 3000.04115391238, 3311.58459987263, 
    3311.58459987263, 3979.36880509946, 4320.5301664678, 4386.73134577807, 
    3450.92445737476, 3387.2978515625, 3114.29823439717, 3319.91227025609, 
    3319.91227025609, 3296.73872939792, 2888.66305192277, 4999.27718787381, 
    5471.29152663441, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5404.15511479684, 5452.66807538873, 
    5382.96681124682, 5283.15201708016, 5310.57509767239, 5333.62167333457, 
    5269.33575085598, 5195.21373027288, 5162.09769261952, 5128.21473027894, 
    4911.24860754849, 4913.79884238439, 4730.27531724015, 5232.46309385286, 
    5178.98494884897, 5072.42778535194, 4999.03758917675, 4954.36884058497, 
    4763.81820209991, 4763.81820209991, 4748.06531686451, 4733.91545038687, 
    4623.45540218693, 4393.97963610732, 4240.69557994528, 3995.09867785864, 
    2257.23869070365, 100, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 1767.65452680899, 
    3450.94386916722, 4099.08342211809, 4542.04209957617, 4658.70442183977, 
    5185.09597584027, 5368.34728967148, 5297.29116828811, 5117.18981914939, 
    5077.80517628447, 5073.66401422322, 5024.35470935058, 5019.13342917579, 
    4864.73560304874, 4493.76773895766, 4741.9841574962, 4779.07571895829, 
    4835.11719233179, 5064.03130877509, 5247.44305328868, 5423.9175575724, 
    5500, 5441.42213961797, 5172.26449589844, 4727.11830654443, 
    4025.51589883286, 4543.37315944438, 4639.60625641078, 4639.60625641078, 
    4706.77428058506, 4579.98418698203, 4419.18185522252, 4046.58283475456, 
    3970.0830688422, 3965.44738694613, 3563.18441136069, 3319.65989088003, 
    3099.57004689856, 2384.05126498444, 2379.80487696549, 2631.091998118, 
    2857.38604258104, 3241.65662565874, 3296.20860487586, 2897.86406664522, 
    2191.85384798669, 3169.03915381896, 3169.03915381896, 3789.1920793858, 
    4446.10272091169, 4954.69552919944, 5132.20975904795, 5126.88599987474, 
    5174.00753617878, 5181.50081930819, 5156.38743763797, 5068.01722726427, 
    4897.14884745373, 4102.15073462906, 3387.2978515625, 3387.2978515625, 
    2848.3449812833, 4194.39150875792, 4367.80335589416, 4367.80335589416, 
    4255.58015659521, 3949.15163543251, 2553.36887574786, 1412.00317480215, 
    1050, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    40, 90, 230, 302.029492921295, 880, 1527.05636830172, 2984.81336064114, 
    3375.52706010849, 3185.52598353397, 2703.59399301473, 2338.39100696543, 
    2338.39100696543, 2050, 2050, 2050, 2530.12487545024, 2650, 2650, 2650, 
    2650, 2377.53463480861, 1478.68884277344, 825.529498400984, 
    825.529498400984, 591.455088506497, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 40, 40, 70, 80, 80, 60, -0, -0, -0, 150, 160, 160, 150, -0, 
    -0, -0, -0, -0, -0, -0, 40, 1805.11386238468, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5442.80550569614, 
    5310.52828175974, 4583.96945020067, 4324.59056741724, 4394.40894395567, 
    4394.74921110733, 4394.74921110733, 4974.54020637722, 5494.27561601341, 
    5500, 5500, 5500, 5500, 5417.19363006544, 5430.31986875038, 
    4857.84218701174, 580.953491210938, 4638.07768174306, 4799.04825178272, 
    4889.15183715636, 4320.5301664678, 4320.5301664678, 3794.51242599055, 
    4036.26023292778, 4199.09759741614, 4281.75661755698, 4281.75661755698, 
    4025.82575601475, 3643.24155977078, 3847.41177834363, 5218.98871699945, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5491.00426830096, 5456.97227002994, 5373.21949995997, 5293.70984150579, 
    5239.10468054799, 5378.51945131971, 5347.74225319146, 5356.24011763662, 
    5363.19042644699, 5235.34106250104, 5185.01114787319, 5215.29869817947, 
    5203.35559322063, 4974.04389558674, 5132.08552765536, 5164.16702391743, 
    5188.82010689767, 4999.03758917675, 5073.7307079104, 4959.6114288778, 
    4763.81820209991, 4763.81820209991, 4748.06531686451, 4621.37345083332, 
    4556.32591736234, 4200.00814375496, 3834.58510807368, 3487.50618583966, 
    714.787507887036, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 2308.16792985951, 
    3597.00415893876, 4177.8523536371, 4326.87322265465, 4498.96293723469, 
    4876.02986313675, 5045.07400978945, 5045.07400978945, 4954.36733914526, 
    4835.31820671808, 5038.62472211453, 5019.13342917579, 4985.95207022574, 
    4811.98705139998, 4663.24343722396, 4937.65596667512, 4903.11830745981, 
    5064.03130877509, 5064.03130877509, 5429.39125609047, 5448.53266996428, 
    5361.1734407743, 5254.30684227774, 3596.51229270179, 5042.58216262182, 
    5022.61001968873, 4838.82748976126, 4501.92960089327, 4647.31783489635, 
    4647.31783489635, 4735.78085169926, 4324.42729360604, 4096.06363330076, 
    3999.60531607989, 3882.4035285368, 3621.54774480036, 3589.23230726111, 
    3182.14005652304, 2964.76866978852, 2418.35455390098, 2242.96423050341, 
    2558.16987958323, 2499.72423865193, 2710.3680145276, 2909.01522845717, 
    3266.00061014864, 3261.73464247464, 3423.07964611221, 3864.57998791957, 
    4210.27572408321, 4596.88901337394, 4657.39721417581, 4822.92312592632, 
    5100.04547990982, 5100.04547990982, 5099.27001845865, 5099.27001845865, 
    4473.21246856368, 3311.62790627474, 2368.73740037927, 2848.3449812833, 
    4194.39150875792, 4367.80335589416, 4367.80335589416, 4382.1049147327, 
    3949.15163543251, 2553.36887574786, 1412.00317480215, 1050, -0, 850, 850, 
    1050, 1550, 1550, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 450, 450, 
    550, 880, 1850, 3108.50367083008, 3473.10911381276, 3473.10911381276, 
    3185.52598353397, 3014.05763238236, 2925.72668652395, 2338.39100696543, 
    1850, 1850, 1850, 1850, 1850, 2385.25320746196, 2385.25320746196, 
    1825.68822485784, 1825.68822485784, 1612.11596988352, 610.032254496868, 
    591.455088506497, 591.455088506497, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 0, 40, 50, 60, 60, 60, -0, -0, -0, 150, 1577.3172313359, 
    1577.3172313359, 1062.38116221179, 384.443307861378, 724.538254469148, 
    724.538254469148, -0, -0, -0, -0, -0, 1280.12060546875, 4586.41729003374, 
    5500, 5357.67809402639, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 4540.86640187244, 3371.05235635047, 
    4394.40894395567, 4575.43759134835, 4575.43759134835, 4642.72668732325, 
    5115.89851485824, 5445.24165093725, 5354.71169227059, 5364.62901686414, 
    5313.24816907319, 5020.11822225192, 5012.20473147889, 5107.85907875854, 
    3554.58592437844, 5461.23653564181, 5287.53170193945, 5171.08162853661, 
    3725.27950085873, 3794.51242599055, 3886.25683791082, 4036.26023292778, 
    5010.93304768313, 5098.28900294808, 4942.78644865268, 5104.65118964055, 
    5031.45901893918, 4742.64691112215, 4808.73165561218, 5239.07446582907, 
    5500, 5441.9554720041, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5430.50546515668, 5317.19671101418, 5379.88443737512, 5312.4773011628, 
    5352.77444485391, 5306.00031364075, 5340.62569144725, 5479.82415999547, 
    5429.3829253267, 5390.82687248007, 5410.41289083118, 5315.4805480418, 
    5268.95726655049, 5343.72425318982, 5118.56695038064, 5116.4992755875, 
    4990.61793966211, 4990.61793966211, 4949.22337197195, 4897.21812943967, 
    4964.43040990988, 4787.71146232265, 4763.81820209991, 4747.46719955911, 
    4564.03539357912, 4442.65818032523, 4011.22240952562, 3568.86805544499, 
    2287.87859204298, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 
    1598.19251473167, 3055.33210941264, 3580.21282443215, 4163.97767699025, 
    4419.18185522252, 4484.2311895319, 4762.67971366811, 5010.05589941394, 
    5026.07386424734, 4934.55336920054, 4975.85030758545, 5015.31848038876, 
    4998.34685918368, 4866.45846798083, 4991.73156998549, 4746.44177412389, 
    4928.22824732896, 5013.3148717531, 5410.26342926127, 5391.75721341355, 
    5302.21630890918, 5446.43893298026, 5277.27047052089, 4783.39645922537, 
    5122.56874484056, 5122.56874484056, 5064.78571620425, 5064.78571620425, 
    4985.71633953154, 5111.95724714297, 4834.69223721202, 4726.70805876281, 
    4398.76499840428, 3933.66494048445, 3933.66494048445, 3852.98954494732, 
    3508.53469657205, 3460.15032893362, 3190.69989687216, 2608.59200057721, 
    2223.9741391726, 2090.48019818458, 2118.32211052611, 2710.3680145276, 
    2909.01522845717, 3330.97321669018, 3261.73464247464, 3306.06697379486, 
    3306.06697379486, 3274.81020530473, 3364.48806972374, 4050.35431431786, 
    4496.25599767688, 4608.21993541452, 4890.0830203557, 5099.27001845865, 
    5099.27001845865, 4473.21246856368, 4239.14739275813, 3427.50491803613, 
    2244.66194242854, 3931.07368305514, 3770.31446807029, 1745.91948155658, 
    3017.89672182075, 3017.89672182075, 1624.55243384499, 1050, 1050, -0, 
    850, 850, 1050, 1550, 1550, 1850, 1850, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 450, 450, 550, 880, 1845.85181778795, 3281.27405648891, 
    3473.10911381276, 3473.10911381276, 3289.08326041317, 2925.72668652395, 
    2925.72668652395, 781.251682912977, 607.460387725857, 750, 750, 
    326.990295410156, 339.844358277883, 339.844358277883, -0, -0, -0, -0, -0, 
    60, 60, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 40, 40, 50, 70, 70, -0, -0, -0, -0, 603.882538860719, 
    1577.3172313359, 1577.3172313359, 1337.64719684552, 1162.31879919297, 
    2645.37781280492, 2559.72670625767, 180, 220, 220, -0, -0, 
    270.610395222517, 1369.12234111374, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5049.48709233688, 
    4764.71212974857, 4631.87823547463, 4575.43759134835, 3750.27618038379, 
    4286.96304348563, 4807.18915363896, 4807.18915363896, 5109.42278824253, 
    5122.32229604241, 5122.32229604241, 5122.32229604241, 4629.66288730002, 
    5294.76231156616, 5500, 5434.29236279282, 5366.54592722785, 
    4176.85837743299, 3543.00211581246, 4652.84309091603, 5068.57808341699, 
    5402.23397993946, 5341.40607562626, 5226.07242949822, 5083.00784111748, 
    5083.00784111748, 4843.3931887481, 5326.76273323926, 5198.86395036404, 
    5088.23823376416, 5044.23576416437, 5500, 5500, 5500, 5500, 5500, 
    5396.31214769665, 5121.95209613894, 5341.93220137921, 5500, 
    5302.00120238791, 5494.80856040252, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5488.12315933627, 5374.08565752741, 5451.87092574895, 
    5372.33181157578, 5318.27207950246, 5312.42051165842, 5264.80894223783, 
    5327.52375293243, 5319.62366789802, 5349.40507394923, 5350.43225543515, 
    5334.09349081337, 5328.35349439123, 5338.07556744501, 5293.30649166929, 
    5118.56695038064, 5064.38204824031, 4944.48920149024, 4955.27321354263, 
    5016.20981705229, 4907.13701588027, 4994.33553672176, 4800.81192932357, 
    4705.46420625728, 4621.04724134577, 4456.88728735412, 4257.60720990837, 
    3966.07838077194, 2617.43391778724, 170, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 40, 350, 2421.58499740675, 3039.31124692158, 3609.09620994828, 
    4108.45241965198, 4224.6572496228, 4607.43418266012, 4821.64422264559, 
    4980.24230239534, 4960.46208555583, 5060.31574185492, 5083.91166649417, 
    5082.72755427854, 5089.85368010845, 5084.11902441707, 4973.94786716961, 
    5123.81206996675, 5166.25510571252, 5276.08374580412, 5367.32196251377, 
    5391.63304289196, 5410.91945988097, 5415.79746590943, 5458.13599427853, 
    5426.61921906657, 5409.36467665049, 5344.50058901456, 5315.26313264302, 
    5197.32300927839, 5252.75821031144, 5169.60444310175, 4643.91228312161, 
    4344.6965686778, 4344.6965686778, 4177.27117659458, 3987.46603224993, 
    3736.77835585752, 3644.5030510187, 3682.00349084782, 3157.38717716642, 
    3112.84347764153, 1424.91349323596, 1877.80583132519, 1762.85367448564, 
    1641.93324799029, 1559.66834925541, 1980.3414620959, 2149.75245247122, 
    2149.75245247122, 1156.25889250163, 1760.09272186612, 3637.42120244608, 
    4092.65848866483, 4092.65848866483, 4254.93425797263, 4459.06073699467, 
    4459.06073699467, 4500.42598564902, 4239.14739275813, 4239.14739275813, 
    3246.73378558247, 4051.46024438803, 5088.5269041007, 5109.81796400207, 
    4078.1536549542, 1478.68884277344, -0, -0, -0, -0, -0, -0, -0, 1550, 
    1550, 1850, 2050, 2050, 2584.03891465366, 2584.03891465366, 
    2759.20661343594, 2771.46419932143, 2739.77891138135, 1850, 1350, 1050, 
    450, 450, -0, -0, 1861.66671768316, 2466.66776221529, 2794.73896659585, 
    3255.35679152863, 3273.14111148246, 2919.2014814502, 253.361404418945, 
    -0, 90, 550, 550, 150, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 0, 40, 40, 40, 70, 70, -0, -0, -0, 299.947582708618, 
    1581.42418499214, 1907.53585334894, 1907.53585334894, 1907.53585334894, 
    1162.31879919297, 2664.85099699065, 2559.72670625767, 1465.9918358999, 
    1465.9918358999, 384.939738642918, -0, -0, 60, 1102.98099102449, 
    3177.92569092766, 5500, 5365.83885293489, 5270.99028669923, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5376.54377768091, 4811.25197570971, 4138.67780951532, 4528.22452754171, 
    5033.29592027491, 5107.46641338799, 5229.017091591, 5412.10727679554, 
    5421.46786389469, 5500, 5500, 5500, 5500, 5500, 5275.56449421238, 
    4443.66678679451, 4628.64736437222, 5207.01531175981, 5488.41380122367, 
    5500, 5500, 5500, 5083.00784111748, 5394.24730134304, 5500, 5500, 
    5460.25469286294, 5470.27865902699, 5301.80369426205, 5082.03481861138, 
    5497.02559270175, 5500, 5500, 5500, 5492.35664560069, 5239.10227564132, 
    5111.71457990612, 5410.30495547833, 5481.57685503835, 5384.6927229193, 
    5337.09473619568, 5466.07778427091, 5287.69902604001, 5243.90953561082, 
    5500, 5500, 5500, 5302.88790697286, 5500, 5395.39769782563, 
    4976.17776159005, 5200.78994016751, 5145.77292429043, 5036.53353093166, 
    5245.34366351458, 5218.70457944923, 5476.09186415092, 5273.20220196002, 
    5303.34850628825, 5242.88829037087, 5258.34640333024, 5235.59755090426, 
    4980.2954163074, 4982.94021376275, 4856.2081030024, 4716.48809744467, 
    4716.48809744467, 4664.53564048247, 4635.58827751501, 4628.9584818942, 
    4569.05492933903, 4566.89303566491, 4564.79719724197, 4353.48939939286, 
    3820.32574750543, 3630.92946361908, 276.864961049193, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 40, 370.154968261719, 2659.38264862153, 
    2835.73762309184, 3090.74178595806, 3462.19595886353, 3900.09318260192, 
    4330.59456382268, 4622.810554932, 4779.07571895829, 5020.75445870074, 
    4639.72850508769, 4840.02249450207, 5124.94883708849, 4667.34325412913, 
    5174.26597922756, 5197.29410643095, 5269.43860427323, 5331.81952402013, 
    5352.89573936724, 5361.79396363088, 5353.22132775751, 5413.78106322914, 
    5409.70920048854, 5492.078972922, 5443.41817057833, 5372.82005027213, 
    5361.84922277613, 5304.35575960383, 5195.66992071839, 5207.34180606951, 
    4650.90657062796, 5087.27756818791, 4946.68021441713, 4835.3429545688, 
    4574.16383399285, 4459.94207842029, 4335.88585029655, 4334.97666192181, 
    3986.63529045442, 3113.45696468855, 2683.8928697654, 2124.28353384322, 
    1530.14401682826, 1582.81609941241, 1668.85081544936, 557.584992504036, 
    1202.16586817197, 1439.78624325437, 2789.54549386887, 3550.53899290818, 
    3873.67527900619, 4176.20239649748, 4401.66837108954, 5007.5393336726, 
    4886.00731841915, 4666.60540426885, 4793.9800304728, 5346.85460644665, 
    5371.85723168386, 5345.10708238118, 4051.46024438803, 4862.5793080226, 
    4816.22739134266, 4078.1536549542, 768.295393786641, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 1850, 2050, 2050, 2622.43913736358, 2584.03891465366, 
    2830.17858331053, 2852.09706852064, 2739.77891138135, 1850, 1350, 
    1268.76743640531, 1219.86869350762, 1292.66416858461, 1409.72581199013, 
    1409.72581199013, 0, 1850, 1865.29432589124, 2564.00238610319, 
    2564.00238610319, 687.448416965143, -0, -0, -0, 410, 410, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 0, 40, 40, -0, 50, 50, -0, -0, -0, 299.947582708618, 
    1581.42418499214, 2128.17192162256, 3014.37518884513, 2945.68599801208, 
    989.372636698672, 989.372636698672, 748.637730982349, 2506.58052745905, 
    2518.06509102109, 1643.78420552745, 623.231301883022, -0, -0, 
    908.577786079993, 2669.61807065125, 5500, 5315.21144959599, 
    5219.39080153592, 5268.46146866994, 5500, 5500, 5407.37531109078, 
    5450.7216827416, 5500, 5500, 5500, 5500, 5500, 5500, 5497.53886213942, 
    5500, 5500, 5312.43416668674, 4936.42368161502, 4836.1200049606, 
    5123.80132744763, 5195.45934611862, 5161.17838014291, 5490.53378729586, 
    5500, 5500, 5500, 5500, 5500, 5066.94767635332, 4649.71690918664, 
    4994.30223028979, 5412.9481062632, 5500, 5500, 5346.92389418097, 
    5225.84165545244, 5347.71674246328, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5473.94381368495, 5500, 5500, 5500, 5500, 5500, 5447.60721527874, 
    5412.80307482045, 5495.71808870876, 5500, 5402.68316348733, 
    5389.06317390542, 5183.20027405752, 5266.49321454198, 5207.88934955842, 
    5284.33322154713, 5075.06786134063, 5433.03169769173, 5414.326361837, 
    5463.7566364326, 5220.99184844207, 4976.17776159005, 4976.17776159005, 
    4899.47669457609, 4763.30603960183, 4541.28899717677, 4897.9370117177, 
    5143.41858983545, 5375.90588329914, 5470.84936743481, 5387.0605565696, 
    5283.14193543836, 5217.17248375551, 4980.2954163074, 4989.13423118173, 
    4958.12124555428, 4716.48809744467, 4739.75965146749, 4544.05465216861, 
    4446.39294677925, 4437.44321081223, 4445.62423409596, 4319.16296011078, 
    4318.4927768179, 4125.68538361722, 3552.18531924069, 2117.34751843701, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 40, 350, 
    1913.24200248399, 2387.14009498566, 2340.39370132507, 2815.31053971462, 
    3498.28073072544, 4036.36273492269, 4036.36273492269, 4639.72850508769, 
    4639.72850508769, 5028.28528168975, 5054.79321645082, 4952.48115133659, 
    5143.41858983545, 5192.16992160785, 5236.07249982981, 5273.57148280206, 
    5274.1804246818, 5249.43991413152, 5262.21228791842, 5292.07564914099, 
    5350.53613011987, 5356.74197996776, 5406.44632142147, 5274.6114783769, 
    5143.41858983545, 4402.70573818403, 4260.8590228139, 4618.8034941342, 
    4650.90657062796, 4889.25934043691, 4985.83837216404, 4829.12129476937, 
    4747.21060530736, 4452.91203839148, 4352.80992925018, 4270.0014508059, 
    4086.3534628009, 3796.2835429095, 3202.47357772414, 2013.6795152968, 
    1524.10942966774, 1582.81609941241, 1582.81609941241, 1657.50197655536, 
    1657.50197655536, 2641.04702665216, 3054.94256249199, 3644.79374030902, 
    3863.92083310841, 4080.29514575055, 4401.66837108954, 5058.58920304941, 
    4867.87069872262, 4666.60540426885, 4793.9800304728, 5159.75546360932, 
    5292.85319076192, 5143.41858983545, 4250.27834514013, 4079.07774156682, 
    4079.07774156682, 3349.04400521109, 402.942120660804, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 495.553629324057, 495.553629324057, 650, 1550, 1850, 
    2808.66018585083, 2848.05298066138, 2400, 1250, 1250, 1632.72145037847, 
    2578.30920183069, 2578.30920183069, 1546.25789094543, 1409.72581199013, 
    0, 1150, 1150, 1150, 833.221376107709, -0, -0, -0, -0, 260, 260, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 782.693477947901, 
    2418.69859717649, 3229.12356137073, 3290.7255144827, 3295.86555058579, 
    2549.42505613294, 2466.66776221529, 2826.94092366, 2826.94092366, 
    2978.4092564626, 1359.10391277954, 40, 40, 1121.77923414952, 
    2171.14041753625, 5500, 5500, 5151.1522329727, 5313.80272145484, 
    5382.89167015676, 5386.27243357935, 5373.9624471111, 5352.2189807718, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5486.26471143345, 5102.90562457836, 5123.80132744763, 5500, 5500, 5500, 
    5500, 5500, 2761.48531639985, 4927.68287286693, 4927.68287286693, 
    4370.49824254822, 5012.38577864191, 5500, 5500, 5500, 5500, 
    5331.82855979701, 5403.59694570381, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5439.76332625033, 5363.34992113622, 
    5423.26897125918, 5500, 5500, 5437.09333741768, 5384.417720333, 
    5274.23306369577, 5212.63844856299, 5267.87690126216, 5376.83857607288, 
    5400.56944960453, 5154.06164964968, 5125.96045844389, 5047.32582429337, 
    4787.33357623623, 4744.5445246852, 4710.54831369341, 4710.54831369341, 
    4649.16410988564, 4604.42242853963, 4634.40210414685, 4672.77236671858, 
    4731.10457537932, 4555.87354394826, 4690.79781441172, 4672.3654865445, 
    4419.18185522252, 4225.20491317775, 4229.14569503725, 4323.89175939117, 
    4312.83055502545, 3959.96072659777, 4003.53541554914, 3846.9806235541, 
    3629.60779216964, 3456.60267593453, 3040.63851545185, 3040.63851545185, 
    2962.34155120925, 2962.34155120925, 2558.86560492922, 550, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 50, 90, 90, 140, 140, 
    425.785466617812, 2388.05438830022, 3800.27626019494, 4439.99525965215, 
    4554.44261634601, 4748.92651424947, 4830.4147003611, 4952.48115133659, 
    5048.22167733199, 5083.87550616628, 5166.38343494461, 5203.10288867419, 
    5160.18700426736, 5121.10558676316, 5200.7362147052, 5209.4964816061, 
    4572.41997132352, 4065.89147763595, 4073.33410400882, 3721.27612304688, 
    3726.68790021752, 4159.94006856668, 4530.22789542051, 4730.06255317601, 
    4789.4622011084, 4947.37781799313, 4971.61111402372, 4781.25304176479, 
    4687.42665269221, 4579.53094441862, 4352.80992925018, 4359.19399030749, 
    4359.19399030749, 3920.67671902433, 3474.29338634069, 2718.05299686344, 
    2220.50553506282, 1973.51337911259, 1894.61889247799, 2299.13594339492, 
    2253.22842819085, 2704.60854424838, 3054.94256249199, 3548.17390562063, 
    3863.92083310841, 4022.85729342828, 4006.63103674706, 4404.36772703333, 
    4693.75012968053, 5113.35421842435, 5113.35421842435, 4899.71255615276, 
    5113.97350881937, 5254.85337307753, 5340.99954793261, 5300.3476456103, 
    4079.07774156682, 3349.04400521109, 928.02522314794, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 40, 350, 1478.68884277344, 2631.72573181078, 
    2760.74151612467, 2794.78195553759, 2605.40963353482, -0, 1250, 
    1632.72145037847, 2578.30920183069, 2578.30920183069, 1546.25789094543, 
    0, -0, -0, 650, 650, -0, -0, -0, -0, -0, 210, 210, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 2418.69859717649, 
    3177.31784759196, 3243.05480048537, 3243.05480048537, 2624.69934803557, 
    3546.22352226187, 3423.84076652799, 3594.14274947404, 3300.17303348703, 
    1411.39339752854, 40, 40, 1204.80827787095, 1241.04603027255, 
    3736.2583354771, 5500, 5500, 5209.98954718568, 5199.50706860803, 
    5280.77999540082, 5238.8436839217, 5253.84185937607, 5329.79884848084, 
    5470.65295715725, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5222.19738159041, 4731.64752924737, 5223.69822293899, 5365.27937785067, 
    5477.32653588348, 5500, 5382.19754659876, 2392.8184540144, 5500, 
    5202.49793796231, 5129.42278239258, 5469.63181166241, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5465.08847615697, 5294.70125536378, 5415.21608022488, 
    5427.38853159314, 5500, 5375.34610381455, 5288.16405469162, 
    5270.60681761282, 4696.44895178471, 5257.20316380099, 5275.37117629753, 
    5282.28564350993, 5194.50429953288, 5125.96045844389, 5022.33559021971, 
    5057.27978573479, 4954.4934559412, 5110.18989840362, 4951.12327809073, 
    5123.68257175295, 4852.40186593518, 4664.21159769676, 4704.7275357794, 
    4703.0225846691, 4589.17933545522, 4533.39354280014, 4445.22039111072, 
    4297.70030896214, 4194.57919244279, 4099.35246362854, 4001.07785590758, 
    3944.25492035913, 3853.62254281299, 3739.2973683011, 3579.98561428294, 
    3455.25033950311, 3223.56465273313, 3107.57190354874, 3154.14952294923, 
    2630.0950131275, 2643.09136179928, 2643.09136179928, 550, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 140, 140, 50, 
    140, 2266.863451998, 3175.33331329546, 3497.21619812172, 
    3897.31723365164, 4440.4727928723, 4641.58152408516, 4837.48618633413, 
    4984.6957231874, 4972.99713307389, 4977.96153711168, 4730.60026757273, 
    4919.04856020589, 4889.48852355269, 4958.62986560659, 4335.61717528916, 
    4041.40151663801, 3174.29635324872, 3432.36288190208, 3903.47237851819, 
    4558.49546877835, 4768.18469648456, 4902.38748684381, 4931.64423719712, 
    4917.15130072564, 4905.25356754764, 4795.45104981751, 4678.20114758192, 
    4476.80444811394, 4340.0214745808, 4359.19399030749, 4399.06665393779, 
    4012.4143292355, 3854.2438971654, 3309.81556918399, 2626.17089832179, 
    2288.08083745065, 1894.61889247799, 2242.66735095028, 2547.78323610602, 
    2873.56017852434, 3317.69107604188, 3548.17390562063, 3735.83694873752, 
    3735.83694873752, 3595.96907035686, 3675.30024756466, 4466.76131756313, 
    5113.35421842435, 5113.35421842435, 4963.99151431876, 5164.8095443174, 
    5330.91422738345, 5347.29511772297, 5249.43607318662, 3065.78548661781, 
    3175.5446543715, 1008.471410908, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 40, 1478.68884277344, 2565.48213236658, 2550, 2683.23341343172, 
    2615.50619077256, 0, 985, 998.018983942509, 998.018983942509, 0, -0, -0, 
    -0, 480, 650, 650, -0, -0, -0, -0, -0, -0, -0, -0, -0, 180, 
    656.90881385992, 656.90881385992, 641.500005998289, -0, -0, -0, -0, 
    240.561416625977, 1450, 1762.59335750926, 1763.50839409499, 
    1454.12072823282, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 425.785466617812, 
    1003.80275890641, 1484.98110495847, 2624.69934803557, 3550.31608409607, 
    3467.5430449472, 3693.20512554389, 3300.17303348703, 2277.75786007126, 
    -0, -0, -0, 60, 1074.81554283494, 2512.95460103342, 4427.24685979802, 
    5500, 5500, 5061.17406184948, 5018.77468813783, 5087.70541714126, 
    5217.10699688685, 5343.44826975707, 5292.96230113963, 5451.90175309996, 
    5481.29516648737, 5486.16184818749, 5448.78062973323, 5500, 5500, 5500, 
    5485.01486470985, 5207.62359403881, 5079.62112516098, 4779.07571895829, 
    5014.80769442128, 4957.61710646844, 5196.67240264642, 5500, 
    2621.42111182486, 5500, 5377.07080006989, 5129.42278239258, 
    5301.50590646636, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5321.81140617512, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5403.89634811281, 5418.44064468193, 5500, 5409.42240480011, 
    5343.7670107254, 5295.58216615451, 5439.67387681021, 5380.41855319955, 
    5335.93793884765, 5419.80576615543, 5270.15190682318, 5185.29786051516, 
    5022.33559021971, 5088.21730853414, 5088.21730853414, 5088.21730853414, 
    4951.12327809073, 4802.51398261262, 4810.16178774669, 4664.21159769676, 
    4420.90451291616, 4554.29173121861, 4459.54291619602, 4329.81907814643, 
    4353.7470749278, 4128.80674283622, 4161.49684410373, 4036.16798145613, 
    4007.51591109129, 3989.11012902597, 3899.61910270725, 3678.94578444491, 
    3496.68899379769, 3606.46355309833, 3371.48874953515, 3197.01659944444, 
    3196.08630333252, 2819.43895627994, 2643.09136179928, 2643.09136179928, 
    315, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    40, 100, 140, 140, 140, 140, 919.053638408483, 1552.27981095526, 
    1872.0268245299, 2780.92176380007, 3531.11429991868, 4270.7173833784, 
    4387.76040364532, 4387.76040364532, 4361.53542257451, 4338.17885366877, 
    4696.50484212836, 4618.21548365607, 3742.24708201151, 2681.38337557688, 
    2143.41355604805, 2762.63296612624, 3281.63703005327, 3903.47237851819, 
    4534.20438248416, 4768.18469648456, 4862.67699852649, 4873.8170039588, 
    4868.57154852796, 4877.33795528503, 4869.51811588893, 4555.13373721637, 
    4246.17366721401, 3762.74248786622, 4108.3507422288, 4137.35282760538, 
    3990.16388312354, 3807.58039888379, 3392.68836842111, 3047.52966600829, 
    2713.27442344581, 2240.77681157926, 2242.66735095028, 2736.90914717819, 
    2873.56017852434, 3317.69107604188, 3556.3438464213, 3535.75227927008, 
    3646.32297703989, 3567.44809198166, 4031.00612776669, 4125.9172908059, 
    4384.63061149358, 4836.57863403192, 4963.99151431876, 5178.91293700599, 
    5354.20441993747, 5299.79542158675, 4442.9324451232, 1603.66521414229, 
    1603.66521414229, 1008.471410908, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 327.909353794418, 1589.84791105535, 2263.76863841736, 
    2615.50619077256, 2725.19413532511, 1415.92336539055, 985, 985, -0, -0, 
    -0, 230, 230, 480, 480, 480, -0, -0, -0, -0, -0, -0, -0, -0, -0, 180, 
    656.90881385992, 1211.28078135842, 1697.12502302956, 2126.90092412782, 
    2096.25319649454, 1939.91402838438, 1917.81264172573, 1922.42002461917, 
    2092.53269301321, 2058.6329902323, 1762.59335750926, 1454.12072823282, 
    -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    1436.52416241863, 3393.95723214103, 3583.13740534935, 3227.26035008689, 
    2277.75786007126, 220, -0, -0, -0, -0, 170, 240.561416625977, 
    2269.91911295663, 5061.17406184948, 5061.17406184948, 5112.67633416182, 
    5112.67633416182, 5150.44404143628, 5263.1802071895, 5409.93340125305, 
    5410.67711867383, 5403.96172200102, 5500, 5496.98348326345, 
    5436.11358175834, 5414.82693438877, 5500, 5500, 5500, 5500, 
    5449.25205727958, 5005.80297400153, 4857.09965663778, 5448.41862995388, 
    5495.57415409859, 3242.74037471342, 5500, 5194.37002676304, 
    5163.12953397217, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5470.16442806743, 5455.12494326077, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5499.83402176945, 
    5383.28548165467, 5381.69373478228, 5433.58688928083, 5360.60144359862, 
    5198.40862332559, 5459.79468020244, 5500, 5400.24153207451, 
    4924.10302099748, 5088.21730853414, 5088.21730853414, 5093.55655021104, 
    5094.65327889478, 5069.85831590953, 4804.48927980577, 4595.52697087017, 
    4605.99835992559, 4384.08158023047, 4379.34633297751, 4311.57197295718, 
    4277.38324567044, 4220.58594445001, 4166.24098671465, 4045.83434317464, 
    4018.5637219194, 3964.4828108735, 3872.55831173916, 3721.27612304688, 
    3609.40132589441, 3495.53885479527, 3371.48874953515, 3255.37242942798, 
    3070.55216686588, 2873.33115917617, 2950.87918800581, 2859.52693075893, 
    355, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 100, 140, 140, 140, 140, 140, 410, 650, 650, 985, 1398.31454972698, 
    2926.96019935289, 3536.6146467915, 3388.38117539175, 3925.9862606599, 
    3875.51552178243, 3282.34891678627, 1866.87403457739, 170, 70, 
    240.561416625977, 2845.74250281978, 3837.58892844316, 4332.01464748275, 
    4459.61732655641, 4760.40093948081, 4662.44891028715, 4812.49744958941, 
    4799.11921821724, 4824.66373757539, 4609.53580266803, 4200.97066188983, 
    3831.67281228223, 3959.54869481899, 3529.67707130922, 3626.85592881992, 
    3660.12189350226, 3570.04418055945, 3268.46320957478, 2883.35842368966, 
    2299.62770002888, 2091.31523331475, 2736.90914717819, 2736.90914717819, 
    3104.36026264958, 3309.34871662521, 2896.9287251521, 2551.16252235306, 
    3703.28325223094, 4198.74788587276, 4212.91371378704, 4212.91371378704, 
    3644.89301390049, 4066.37981347831, 4965.73371510261, 4866.65048910806, 
    4646.91808412633, 4442.9324451232, 4233.49870893579, 4241.08205965444, 
    1205.3730875484, 485, 485, 485, 485, 485, 230, 230, -0, -0, -0, -0, -0, 
    -0, 0, -0, 1450, 1415.92336539055, 1415.92336539055, 315, -0, -0, -0, -0, 
    230, 230, 480, 480, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    561.393870373234, 1211.28078135842, 1697.12502302956, 2033.51331957481, 
    2118.87790053842, 2160.12061116943, 1917.81264172573, 1922.42002461917, 
    2106.74400796201, 2038.29149311131, 753.47203223552, -0, -0, -0, -0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 608.204723139333, 2163.84062722417, 2090.96749967482, 
    1068.77367355403, 220, 70, -0, 80, 1086.15579679338, 1086.15579679338, 
    270.610395222517, 180, 402.898573978307, 3914.2542323696, 
    5112.67633416182, 5112.67633416182, 5500, 5228.71205872617, 
    5102.89607788252, 5143.41858983545, 5272.98659105091, 5303.52445318286, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5434.21537014364, 3242.74037471342, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5481.69722190124, 5373.79239046475, 
    5416.25593299475, 5346.47338722845, 5301.46380415743, 5254.90386899421, 
    5248.31412131023, 5318.54206793468, 5297.61158064131, 5296.24429444773, 
    5381.89096523999, 5370.95430836386, 5261.67473707582, 5209.09561254307, 
    5259.77030537539, 5260.58403665714, 5173.92670943071, 5103.36682955807, 
    5000.12260410043, 4974.48453856889, 4856.55027952399, 4613.85220426378, 
    4618.34174227993, 4343.07872631123, 4267.83990808051, 4385.86191207411, 
    4193.92139110942, 4184.32253932863, 4131.90200272625, 3990.97784040899, 
    3970.59749310972, 3819.39934230187, 3767.06724870925, 3681.53410850866, 
    3576.06470266782, 2599.6739553561, 2676.49796489373, 2776.00856660753, 
    2890.93953921779, 2915.96895004784, 2825.33440682898, 355, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 
    40, -0, -0, 40, 70, 70, 210, 210, 210, 294.462890625, 1355.37800617976, 
    1948.12288578358, 1948.12288578358, 461.816626598226, 110, 80, 60, 60, 
    2726.04792045947, 3726.65982904536, 3786.16198213809, 4137.03733216239, 
    4674.75644896692, 4691.31273161807, 4767.16703098079, 4767.16703098079, 
    3683.1781633273, 3826.0181017275, 4109.00300726629, 4144.12288098328, 
    4018.12646489169, 3813.62033990039, 3445.21548499598, 3513.66927872397, 
    3489.46627742243, 3173.72020129554, 2789.89461572067, 2691.13581257075, 
    2267.39269533808, 2438.25371562671, 2747.26281414698, 2747.26281414698, 
    2894.03202538836, 3364.79029075215, 3238.90532098892, 3703.28325223094, 
    4122.85504208618, 4396.5156316856, 4396.5156316856, 4396.5156316856, 
    4065.89147763595, 4866.65048910806, 4916.34790657649, 4422.19448270919, 
    4392.87075967718, 4392.87075967718, 4233.49870893579, 4108.07937153275, 
    4108.07937153275, 4800.07730073825, 4880.96930169055, 4649.22300843847, 
    4234.27454674361, 1723.22878906739, 230, 40, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 50, 90, 506.495873342338, 506.495873342338, 220, 
    1024.98282624745, 1024.98282624745, 997.028238330557, 997.028238330557, 
    -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 378.684052958572, 1068.77367355403, 1068.77367355403, 
    471.320821889931, 80, 0, 80, 1161.28758740964, 3065.78548661781, 
    3120.6099643616, 2725, 341.90213998116, 253.361404418945, 
    459.451469285212, 2681.40271423809, 5500, 5500, 5098.03243678519, 
    4932.61413111386, 4996.34094423389, 4877.26339424593, 4796.02344296714, 
    5192.51549961194, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5307.29813490472, 5295.77898223321, 5394.44581038476, 5227.26760608547, 
    5174.92489185305, 5143.57544501159, 5104.63941351433, 5148.92466793955, 
    5171.01212100176, 5223.63334191327, 5215.33760551089, 5207.83228873618, 
    5202.56263441903, 5241.94578142287, 5215.76031008735, 5248.7926689276, 
    5192.08128771331, 5192.74761953363, 5158.42183086641, 5118.99910793774, 
    4963.41780142748, 4817.43031669686, 4795.66568010002, 4670.26435005172, 
    4621.1119192065, 4571.74343494587, 4469.13685271863, 4357.01802127588, 
    4355.5180331329, 4304.97584174874, 4219.86824211648, 4223.31216406661, 
    4133.00891795456, 4004.31608836766, 3800.29914264068, 3556.73278994791, 
    3084.51290696571, 2533.71627957903, 2642.53846225864, 2804.36325363461, 
    2879.2900239536, 2733.97340475125, 2268.34782201321, 355, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 210, 210, 210, 210, 210, 100, 90, 80, 80, 80, 80, 70, 
    587.140122884625, 2191.85384798669, 3001.08758011801, 3721.27612304688, 
    4563.23365184907, 4725.02094236772, 4691.31273161807, 4659.9517666989, 
    4614.18846805776, 4437.84874775814, 4491.63179884038, 4321.97224459562, 
    4403.80090722506, 4163.08815308037, 4065.89147763595, 3743.18871455568, 
    3691.11979872939, 3268.36624527129, 3105.18118925007, 2924.46864509118, 
    2303.80711892699, 2194.57252445333, 2937.29133108035, 3000.55227014129, 
    3040.0177888873, 3315.89969326733, 3799.7418203521, 3928.43990631137, 
    4345.2439374107, 4396.5156316856, 4396.5156316856, 4396.5156316856, 
    3906.82853690828, 4663.32838396905, 4600.65351422648, 4615.25847772487, 
    4392.87075967718, 4392.87075967718, 3670.93620832819, 4765.57123067861, 
    4765.57123067861, 4951.21583137741, 4895.28050535877, 4604.24985398189, 
    4234.27454674361, 1723.22878906739, 120, 40, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 40, 40, 40, -0, -0, 0, -0, 0, -0, -0, -0, -0, -0, 
    -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 542.614650548053, 542.614650548053, 506.413097905128, 200, 0, 
    40, 1720.84480296144, 3253.25149184514, 3302.62206577075, 
    3306.36900576271, 3371.73664950956, 3258.67933297975, 2725, 480, 
    2518.78488077372, 4419.18185522252, 4932.61413111386, 5094.3355719826, 
    4917.97286048464, 4736.63963412132, 4949.72774227191, 5143.41858983545, 
    5409.86879812733, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    2810.51717508525, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5450.63333470365, 5500, 5500, 5500, 5500, 5500, 5500, 
    5390.63861317858, 5500, 5500, 5500, 5500, 5486.18357628058, 
    5383.42468167104, 5338.59453489314, 5215.01580978446, 5121.01348512029, 
    5011.3963897027, 4998.2494720351, 5006.51446941282, 5077.54303974094, 
    5124.39822356124, 5128.53311459267, 5128.53311459267, 5288.56810608923, 
    5246.73787084855, 5232.94043020738, 5272.82468767709, 5202.2097843245, 
    5170.84497123772, 5029.23282512662, 5035.42254976318, 4963.36287886639, 
    4832.27913255505, 4802.2609156317, 4721.51731551426, 4587.35869738783, 
    4496.70168807873, 4444.04588221801, 4369.50540918674, 4298.78055029206, 
    4249.11701807405, 4226.17183057213, 4192.79598374401, 4109.25299084766, 
    3909.21755530012, 3829.28534456476, 3395.17322438906, 2711.46195934008, 
    2317.28462055921, 2525.67069025481, 2728.61685818447, 2728.61685818447, 
    2659.9114617034, 1983.9441789969, 150, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 
    40, 130, 140, 150, 150, 90, 90, 90, 60, 100, 100, 90, 80, 100, 1150, 
    1150, 985, 1341.34845729854, 3770.2484327786, 4011.8355933077, 
    4450.51159137726, 4513.75724632954, 4646.80172448333, 4530.61415341145, 
    4580.02248620154, 4390.30789360063, 4227.23928399928, 4132.86135939777, 
    4100.66945985931, 3905.59590273844, 3553.7160975538, 3330.21403226727, 
    3205.78943979219, 3041.14131020629, 2645.57211838466, 2792.11079429091, 
    3076.29922723107, 3220.95389236629, 3770.88966508943, 4009.96624308098, 
    4222.32022960908, 4653.43458957793, 4617.42481915019, 4144.6084295607, 
    4247.04741600706, 4482.08429377265, 4493.09841074183, 4613.58256359772, 
    4613.58256359772, 4147.23667723678, 4269.24608430867, 4269.24608430867, 
    4765.57123067861, 4765.57123067861, 4760.29175259183, 4705.35100215565, 
    3891.58792054794, 446.137172106597, 140, 60, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, -0, -0, -0, -0, 
    -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 506.413097905128, 506.413097905128, 374.502888602588, -0, 
    314.274068783434, 1720.84480296144, 1833.00053044869, 3042.76564565658, 
    3295.51777030009, 3302.95765593392, 3349.66633126752, 2725, 2725, 2725, 
    2725, 2731.19947353971, 4917.97286048464, 5011.76112466895, 
    4880.3301499577, 5104.52122604408, 5204.42177430385, 5208.63030334165, 
    5431.94078337637, 5500, 5500, 5500, 5500, 5500, 5500, 5443.11413407775, 
    3160.63875669116, 5500, 5500, 5500, 5389.54149217261, 5500, 
    5399.09005471129, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 5500, 
    5500, 5500, 5355.9133924136, 5500, 5401.81757007084, 5472.66949528761, 
    5398.87261699386, 5327.95266616781, 5338.14699398579, 5267.56262707998, 
    5152.02678284221, 5072.10007327849, 5112.75755698322, 4935.11764818943, 
    5015.57033362158, 4976.27803329774, 4990.32125172537, 5029.4219626644, 
    5046.12914600433, 5152.26130483332, 5143.41858983545, 5148.34304336728, 
    5185.8691367317, 4884.93633990805, 4910.54866520841, 5016.2568146497, 
    4956.21230709856, 4832.55724934394, 4822.02926854784, 4740.40535198044, 
    4624.12605076301, 4419.18185522252, 4456.33643176637, 4386.41361717062, 
    4301.51176650271, 4226.708381579, 4142.62469952496, 4102.81370982587, 
    4095.67441722416, 3853.38158133828, 3928.23623990325, 3616.50679727179, 
    3131.00434082432, 2844.65957688961, 2799.64284394603, 2661.25930368276, 
    2694.55211092767, 2647.55869762882, 2385.19372013677, 1280.12060546875, 
    50, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 60, 60, 130, 130, 130, 130, 130, 80, 40, -0, 
    -0, 130, 130, 130, 110, 180, 1150, 1150, 985, 253.361404418945, 
    1825.85730792728, 3790.92593386481, 4241.51509277024, 4652.67580349765, 
    4623.23334190601, 4546.36939558212, 4487.02500516891, 4301.86341085367, 
    4311.56447355868, 4129.37283723845, 4108.59594824824, 3930.25274390503, 
    3707.03766335583, 3501.59865629912, 3269.98117933012, 3036.50564152828, 
    2645.57211838466, 2676.80476871288, 3280.76880870975, 3555.27839220712, 
    3878.11129304954, 4358.23463935475, 4222.32022960908, 4427.78384018727, 
    4529.41854697929, 4306.74992937606, 4292.28728312564, 4630.44239615523, 
    4685.99164189565, 4749.27222938507, 4664.3805109057, 4147.23667723678, 
    4269.24608430867, 4269.24608430867, 4344.47182381346, 2778.00548636967, 
    2299.03354037694, 964.941070857491, 150, 120, 60, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 374.502888602588, 374.502888602588, -0, 
    314.274068783434, 402.778911781622, 667.797503219974, 1101.54602050781, 
    2025, 2025, 2725, 2725, 2725, 2725, 2725, 2725, 2725, 4880.3301499577, 
    4885.08225706819, 5104.52122604408, 5500, 5498.57280906161, 5500, 5500, 
    5500, 5500, 5500, 5500, 5469.49242762431, 4596.8600746544, 
    4688.13453798461, 4944.31795426481, 4944.31795426481, 4439.48391003288, 
    5076.86858656907, 4867.87542569876, 4919.17344165886, 5344.89729460328, 
    5489.29832915564, 5433.23745586902, 5390.33974058927, 5383.58795192883, 
    5362.97198204687, 5396.26161138439, 5353.33168323296, 5477.3183896756, 
    5445.12193053414, 5445.88215091488, 5143.41858983545, 5216.05087861862, 
    5326.31229422084, 5227.50683234761, 5432.20001714591, 5394.63087749597, 
    5249.83817266423, 5168.9996720473, 5038.29458642829, 4934.28368903323, 
    5012.50336487478, 5003.16832559398, 4874.88931199369, 4938.10324810739, 
    4981.45883942459, 5066.8790805856, 5010.23450146119, 4926.61026664442, 
    5018.66137502585, 5024.64634810032, 5068.62218276609, 4906.08915032492, 
    4779.07571895829, 4832.69585696114, 4740.09363287904, 4670.63365833516, 
    4628.70611874629, 4472.61291741454, 4361.68133245924, 4276.18936372625, 
    4290.56604753172, 4262.18725533432, 4161.20507269766, 4008.70425960392, 
    3969.17016261376, 3969.17016261376, 3949.85477609866, 3988.33088668106, 
    3785.02013424849, 3450.79981268958, 3236.67540183724, 3025.69793014461, 
    2834.58838008121, 2514.09743892368, 2492.77244297399, 2595.02475079746, 
    1321.56743967994, 130, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 0, -0, -0, -0, -0, 60, 60, 130, 130, 130, 
    -0, -0, -0, -0, -0, -0, 200, 200, 190, 609.556179526824, 
    1665.28137658092, 1964.79781461131, 1964.79781461131, 985, 
    1204.22927289781, 3140.3800218576, 3972.67448674589, 4399.77254894988, 
    4472.80646454617, 4488.10232407733, 4549.69020856287, 4367.07276664145, 
    4301.86341085367, 4310.50358856938, 4309.53038588538, 4218.55603722854, 
    3974.89546409646, 3707.03766335583, 3569.10877201131, 3269.98117933012, 
    2616.62908274686, 2239.72942145397, 3135.09151752944, 3418.64362984148, 
    3690.79257489703, 3983.97942628006, 4141.31744025697, 4221.31316349781, 
    4221.67883750448, 4306.74992937606, 4400.68807055719, 4292.28728312564, 
    4749.42688831938, 4749.42688831938, 4685.99164189565, 4420.56482862251, 
    2570.8151028522, 2570.8151028522, 1672.08023690913, 298.454233597761, 
    150, 150, 140, 130, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 220, 220, -0, -0, 150, 428.093183033817, 
    868.328270522663, 1650, 1650, 1850, 2025, 2025, 2025, 2725, 2725, 2725, 
    2725, 1650, 1650, 5500, 5435.86780476046, 5419.7643271038, 
    5416.51635455947, 5473.60715825733, 5500, 5500, 5430.72258614663, 
    5077.66979407893, 4292.90755988422, 4688.13453798461, 5033.3290373586, 
    4944.31795426481, 4655.41206534547, 4911.96740422289, 4847.11304951316, 
    4891.76343647179, 4891.76343647179, 4887.6248476582, 4800.45745378672, 
    4878.47263417037, 4939.50520266624, 4733.62605065618, 4986.47731477266, 
    4850.87764276152, 5025.7019493705, 5064.71427040648, 5067.22109285618, 
    5104.07339876271, 5104.07339876271, 5185.97129877299, 5315.86686358809, 
    5290.29972172185, 5318.28941364392, 5228.80449594566, 5117.22284158262, 
    4956.24292966067, 4876.07085357525, 4914.69204698654, 5021.08642984908, 
    4862.69675210239, 4832.94729572495, 4915.28916717636, 4846.95592202879, 
    4899.99495344857, 4899.54764187765, 4887.42518079947, 4940.55426701545, 
    4911.42259992136, 4751.34403568143, 4751.34403568143, 4717.26223879102, 
    4699.07505863334, 4609.22044026244, 4370.5666238126, 4272.45996783422, 
    4186.76770976835, 4149.25815050684, 3905.94508832012, 4022.25559130007, 
    4049.3365525545, 3864.90528726933, 3913.84822308725, 3909.24446563776, 
    3758.68910359282, 3539.83272045638, 3652.7563204934, 3311.26797894586, 
    3044.02879432246, 3025.69793014461, 2496.42676755383, 2363.65217696896, 
    2326.81278255333, 1046.32314316786, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    60, 60, 130, 130, 130, 40, -0, -0, 0, 0, 100, 254.743272125118, 
    274.691451248024, 326.990295410156, 1283.50280208666, 2180.45025285735, 
    2180.45025285735, 1964.79781461131, 3175.70360722713, 3479.73396518531, 
    4083.92075140881, 4352.12773673655, 4376.98423585481, 4376.98423585481, 
    4232.49722997329, 4228.87467830104, 4216.95369770823, 4133.16191125856, 
    4005.54726632682, 4043.35882946069, 4043.35882946069, 3697.18159288423, 
    3680.70812888649, 3277.10293148083, 3143.19218518745, 2954.27348361819, 
    2799.45500696531, 3388.6312412044, 3695.44546697962, 3836.68170030435, 
    3983.97942628006, 3990.68479554499, 3980.80167918311, 4039.35667411646, 
    4259.59820802088, 4231.39460544567, 4686.64538211992, 4749.42688831938, 
    4760.800439949, 4405.63367276954, 3053.35337847641, 1445.97742602243, 
    614.009871877704, 110, 140, 140, 140, 100, 90, -0, -0, 0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 474.262316119944, 568.243402734782, 
    896.273136133496, 1350, 1350, 1350, 1350, 1350, 1350, 1350, 
    508.704911204077, 357.586429963496, 40, 429.718746352964, 1650, 5500, 
    5500, 5348.96625485535, 5491.47351533559, 5500, 5500, 5159.01994769565, 
    5015.27603884895, 3084.40438875502, 4209.4951811828, 4498.12845138932, 
    4551.47925199788, 4492.95093885319, 5120.63789058113, 4781.46895357338, 
    4407.60247949866, 4906.62603246718, 4891.76343647179, 4887.6248476582, 
    4800.45745378672, 4878.47263417037, 4878.47263417037, 4733.62605065618, 
    4850.87764276152, 4850.87764276152, 5025.7019493705, 5064.71427040648, 
    5067.22109285618, 5104.07339876271, 5104.07339876271, 5111.7701931715, 
    5111.7701931715, 4959.10806235354, 4997.68646806253, 5001.18667106588, 
    4935.8747168675, 4748.73071791598, 4756.14011072862, 4863.38608219863, 
    4844.92358222379, 4789.53856990702, 4899.96318721125, 4851.07758301237, 
    4819.1302287303, 4812.32073453621, 4726.36585718189, 4735.56555238034, 
    4884.30266616793, 4907.18020404357, 4751.34403568143, 4751.34403568143, 
    4687.69608057563, 4606.09621933566, 4447.830287701, 4369.13323598012, 
    4249.11974727418, 4127.98600026065, 3877.42353952686, 3268.71646207341, 
    3281.24730676432, 3931.24824782918, 3741.36786411583, 3678.22305565882, 
    3659.40203966272, 3659.40203966272, 3697.44220187893, 3501.89418741219, 
    3281.70057789029, 3027.23477218443, 2794.69571876551, 2124.5787953193, 
    1924.42352743064, 558.622626355185, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 40, 40, 40, -0, -0, 50, 230, 254.743272125118, 
    254.743272125118, 274.691451248024, 392.524633296121, 1566.65627015718, 
    2451.30853440563, 2451.30853440563, 1917.2620092025, 3899.32625160607, 
    4183.75314113791, 4312.84813985528, 4352.12773673655, 4393.47252143148, 
    4312.82693551439, 4150.93242134329, 4103.47671969883, 3740.46003154601, 
    3500, 3500, 3500, 3500, 3500, 3500, 3500, 3500, 3500, 3500, 
    3650.90222930478, 3844.53154300782, 3938.47926401987, 3854.10200865649, 
    3732.38770642085, 3621.97694691315, 4038.18552248789, 4038.18552248789, 
    4656.72124246813, 4741.36885335198, 4686.64538211992, 4258.71339345375, 
    2662.46938615504, 2667.27704891992, 1445.97742602243, 614.009871877704, 
    130, 120, 120, 110, 100, 60, -0, -0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 60, 628.944454018296, 1112.70482593524, 
    1301.45385087648, 1312.31356529619, 1255.99337442069, 1167.69955155953, 
    1141.63718031219, 1013.91526608731, 922.099158431217, 655.601240161705, 
    508.704911204077, 357.586429963496, 40, -0, 521.60970891522, 
    3122.68409518234, 5500, 5500, 5450.31168700234, 5300.34246433514, 
    5296.18358949754, 5039.44294539632, 4082.77764971119, 2490.03518691714, 
    3721.27612304688, 4075.19484255245, 4298.62385644702, 4298.62385644702, 
    4781.46895357338, 4781.46895357338, 4407.60247949866, 2481.77543899958, 
    2481.77543899958, 2207.97012589542, 586.037685571596, 220, 1050, 1050, 
    170, 170, 140, 3886.95793966352, 4282.69922572992, 4095.58050891964, 
    4373.98991487441, 4969.62202763551, 4969.62202763551, 4959.10806235354, 
    4959.10806235354, 4857.24563313677, 4794.85053900844, 4779.07571895829, 
    4719.86200888097, 4594.63069500334, 4620.72162170319, 4468.61666084061, 
    4711.68916731096, 4766.5621538955, 4750.14794054604, 4728.26246360743, 
    4709.58988304788, 4627.00615965341, 4516.69506992784, 4715.2280712742, 
    4709.05354251617, 4730.62053209142, 4704.41733404835, 4532.28376145886, 
    4341.0207370584, 4307.07628577449, 4237.18112820689, 4065.89147763595, 
    3611.61906989787, 3669.29829650224, 3669.29829650224, 3625.17207481451, 
    3656.61014698572, 3645.53778245224, 3617.7358891319, 3621.51453083955, 
    3556.20139015543, 3329.55429345088, 3045.99064877836, 2758.41088867188, 
    2304.56886191035, 1230.16573927958, 160, 140, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 50, 230, 270.610395222517, 
    270.610395222517, 339.927470043108, 1250, 2449.54549020039, 
    3272.65615777736, 3673.88073175881, 3637.279309389, 4118.1509969206, 
    4157.9163196851, 4254.50594136961, 4122.28781658628, 4144.36113777239, 
    4047.88907172642, 3600, 3620.34164622256, 3671.54264504936, 3500, 3500, 
    3500, 3500, 3500, 3500, 3500, 3500, 3500, 3500, 3609.34757125399, 
    3753.51704626204, 3736.20333421387, 3607.72139376148, 3230.21892586132, 
    2821.46655985127, 4023.83643342612, 4023.83643342612, 4681.0533676165, 
    4616.99835481822, 4545.74848153122, 3530.32578322992, 473.92487937901, 
    862.950276135638, 862.950276135638, 408.056682178012, 130, -0, 70, 80, 
    80, 60, 50, -0, -0, -0, -0, -0, -0, 40, 40, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 60, 598.734202044325, 1386.93743337728, 
    1386.93743337728, 1280.12060546875, 1142.91370575806, 1072.15492724578, 
    1076.16149168116, 1050, 1050, 1050, 350.449976032342, 297.499927401743, 
    0, -0, -0, 1920.2645481339, 2493.81184540184, 5500, 5500, 
    5187.35242320704, 4419.18185522252, 3355.72956108196, 3942.52631117457, 
    4419.18185522252, 4574.97851652807, 4075.19484255245, 4220.71661634757, 
    4220.71661634757, 1150, 394.091721755884, 230, 260, 650, 650, 260, 
    1052.57370326329, 1188.64303812999, 3547.83204719149, 3582.84838251418, 
    3519.34565779216, 3177.28383596865, 415, 415, 210, 140, 90, 70, 
    2810.16166888704, 3741.95279290812, 4722.45568223054, 4779.07571895829, 
    4779.07571895829, 4719.86200888097, 4594.63069500334, 4646.3025338435, 
    4498.66188973939, 4623.22610809631, 4667.52287460589, 4603.72273222741, 
    4492.34675268349, 4438.84522164394, 4512.28254137967, 4520.06055750239, 
    4396.23713599182, 3904.37468750071, 3812.82454944023, 3812.82454944023, 
    3702.19402299222, 4160.48027566201, 4192.90685593214, 4152.16382056065, 
    3870.03496564428, 3857.02212595849, 3847.99047035822, 3770.31744065479, 
    3673.68896658216, 3695.3843702006, 3551.91252599736, 3549.16901947505, 
    3493.74562897578, 3459.21571190035, 2962.08135266663, 2700.26830745778, 
    2466.66776221529, 355, 110, 110, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 120, 210, 270.610395222517, 
    270.610395222517, 1250, 2386.1225307933, 3317.56456013077, 
    3723.13650067864, 3911.3073119496, 4035.58771505973, 4066.73734704634, 
    4089.33322822243, 4075.74423049284, 3981.12658930034, 3500, 3500, 
    3586.56711498155, 3708.61663428952, 3710.22237325444, 3500, 3500, 3500, 
    3500, 3500, 3500, 3500, 3500, 3500, 3500, 3603.44357466989, 
    3603.44357466989, 3572.41264395609, 3737.89690023388, 3737.89690023388, 
    3495.58758033645, 3347.54405021062, 3262.7035520751, 3956.91278228112, 
    3956.91278228112, 3568.20365552467, 2698.61230600042, 2575, 
    359.14954922941, 359.14954922941, 150, 70, -0, -0, -0, 50, 50, 50, -0, 
    -0, -0, -0, -0, -0, 40, 40, 40, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 40, 40, 50, 1075.29918161392, 1386.93743337728, 
    1386.93743337728, 1375.52242409778, 1142.91370575806, 1072.15492724578, 
    1050, 1050, 1050, 1050, 140, 140, -0, -0, -0, -0, 1478.68884277344, 
    3801.86568222254, 4187.47787676683, 4187.47787676683, 3105.32845952125, 
    3355.72956108196, 3942.52631117457, 4419.18185522252, 4548.23332191218, 
    3275, 1650, 1650, 3788.1330045182, 3904.90033567871, 3694.66662071324, 
    3387.2978515625, 2506.67379169443, 2506.67379169443, 1841.2790896279, 
    1052.57370326329, 1445.60147322239, 3828.15157805858, 3837.41130622737, 
    3786.41551337354, 3706.35196651336, 3673.09831850412, 3546.07947037006, 
    3169.86119491424, 2693.5968358049, 1970.25017630914, 1806.60114972507, 0, 
    110, 110, 40, 2132.10002291154, 3042.27385441596, 4160.29696590157, 
    4498.66188973939, 4498.66188973939, 4623.22610809631, 4623.22610809631, 
    4682.4857316339, 4606.82399080195, 4447.51143068066, 4440.32137699062, 
    4577.9109329241, 4396.23713599182, 4161.20181373414, 3812.82454944023, 
    3812.82454944023, 3702.19402299222, 4076.76998729136, 4109.60191770157, 
    4010.48613700149, 3238.83421823148, 3744.75680887058, 3871.8964538492, 
    3825.50203641806, 3617.68428769623, 3532.1652051537, 3392.96618928235, 
    3334.28199481784, 2844.07711767033, 2486.05300373583, 2486.05300373583, 
    1808.17163418686, 475, 110, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 140, 210, 242.20285614065, 1250, 
    2423.87521406058, 3282.88804765196, 3672.44096337103, 3825.55155132253, 
    3906.79895855481, 3848.80965590129, 3500, 3500, 3500, 3518.87097310158, 
    3376.18593536035, 3000, 3000, 2964.99250555538, 2900, 2900, 2900, 2900, 
    2900, 2900, 2980.23573380403, 3161.8580329814, 3245.80390867363, 
    3357.66726217617, 3545.61965265651, 3631.21461222459, 3612.68067729062, 
    3441.19699836255, 3738.72613275517, 3997.63081803751, 3495.58758033645, 
    2424.69716071351, 2407.21016227146, 2431.56024408156, 2508.84485908921, 
    2698.61230600042, 2698.61230600042, 2575, 1550, 1550, 210, 100, -0, -0, 
    -0, -0, 40, 40, -0, -0, -0, -0, 40, 40, 40, 40, 40, 40, 40, -0, 0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 60, 60, 140, 160, 230, 230, 338.078792847833, 1075.29918161392, 
    1391.9757878745, 1280.12060546875, 1050, 1050, 980, 550, 550, 550, 550, 
    301.892217410204, 140, -0, -0, -0, -0, -0, 308.886556165727, 
    2806.39632247483, 3831.05214551185, 3831.05214551185, 3105.32845952125, 
    170, 230, 315, 777, 3475, 3879.73611861882, 3885.576080846, 
    3895.81525007582, 3694.66662071324, 3387.2978515625, 3250, 
    2660.38150701855, 1841.2790896279, 1450, 3816.21639950832, 
    3803.56410727766, 3793.86035586592, 3752.95929997971, 3706.35196651336, 
    3647.38076450992, 3611.68002584289, 3534.32127846786, 3238.23049451872, 
    1970.25017630914, 1970.25017630914, 925.1455676805, 150, 130, 120, -0, 0, 
    70, 100, 140, 434.494506647558, 1198.97913695625, 2486.1673222023, 
    4538.26969149153, 4447.51143068066, 4440.32137699062, 4296.50732689654, 
    4271.48929105142, 4161.20181373414, 2322.67858725228, 3139.50131859953, 
    3695.99190501189, 4012.40335111996, 4012.40335111996, 4010.48613700149, 
    4033.32553183641, 3928.61981326814, 3764.31583852905, 3721.27612304688, 
    3514.52239229933, 3268.63498248386, 3111.8787853092, 3028.33660020028, 
    2893.27519703144, 2486.05300373583, 2203.1243669986, 277.839574916341, 
    277.839574916341, 110, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 50, 50, 50, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 0, 230, 230, 1250, 1250, 2013.62237733191, 
    2846.34957935704, 3342.68493046187, 3626.84555439666, 3626.84555439666, 
    3617.05895893861, 3361.41654327778, 3375.77682243969, 3544.94215348984, 
    3425.90035251464, 3307.62623579888, 3307.62623579888, 3000, 
    2834.72959193745, 2864.34691271083, 2728.78833430566, 2418.6486356974, 
    1898.08297599939, 2008.74985543514, 2483.26772164059, 2710.19521146153, 
    2772.8995693866, 2998.75040465623, 2998.75040465623, 2914.85727196622, 
    2914.85727196622, 2900, 2482.51214287092, 2982.95481937729, 
    3242.2173984491, 3242.2173984491, 3141.57279700325, 2424.69716071351, 
    1329.58021375734, 1425.97477733209, 1906.26191246785, 2575, 2575, 2575, 
    2733.6222650195, 2733.6222650195, 1836.00268145692, 270.610395222517, 70, 
    -0, -0, -0, 40, 40, -0, -0, -0, 40, 40, 40, 40, 50, 50, 50, 50, 40, -0, 
    -0, 40, 40, 40, 40, 40, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 60, 160, 200, 210, 230, 230, 338.078792847833, 338.078792847833, 
    350.789425943846, 336.574096430457, 336.574096430457, 326.990295410156, 
    315, 315, 315, 403.762466065914, 403.762466065914, 301.892217410204, 90, 
    -0, -0, -0, -0, -0, -0, 2807.79690499006, 3831.05214551185, 
    3831.05214551185, 415, 2583.87328747608, 3475, 3570.968181961, 
    3570.968181961, 3475, 3776.01649296945, 3847.10261709723, 
    3868.00416295905, 3859.47870614967, 3858.08423969093, 3846.50099517532, 
    3753.7394186817, 3861.1585435174, 3822.36172864831, 3821.2903340493, 
    3790.60214261742, 3762.37371426658, 3772.52250029416, 3695.27597625236, 
    3599.62419656555, 3460.41328151743, 3394.20145739487, 3238.23049451872, 
    1970.25017630914, 1970.25017630914, 925.1455676805, 150, 130, 120, 80, 
    70, -0, -0, -0, 100, 100, 80, 190, 725.967791892689, 1480.00871507901, 
    4401.92139721904, 4271.48929105142, 4161.20181373414, 4299.28965472685, 
    4299.28965472685, 4275.64048815045, 4041.92117523405, 4012.40335111996, 
    3996.70113182338, 3975.46004794242, 3849.59309804176, 3620.82796835978, 
    3509.62108697159, 3445.97048708414, 3313.38136222851, 3065.78548661781, 
    2796.87176499048, 2802.88128911805, 2269.05472055291, 257.591506312474, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 50, 50, 40, 90, 90, 
    50, 50, 50, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 80, 170, 170, 1127.44248940889, 1847.38975976044, 
    2414.91876681918, 2856.71693634815, 3231.56933744833, 3321.17325635677, 
    3496.19551668933, 3674.41917819842, 3696.98363607819, 3466.05228077865, 
    3182.47995995106, 3356.14769658321, 3355.18409166942, 3328.06337800628, 
    3319.04233238735, 3261.67001797096, 3000, 2967.3409993646, 
    2982.75810803134, 2572.16857180529, 2278.39465179556, 2250, 2250, 
    2309.28900374485, 2435.47179180075, 2671.09156185418, 2868.54007708541, 
    3043.72020971397, 2909.64126824239, 2906.96542249932, 2906.96542249932, 
    2872.01085829926, 2728.7540537158, 2337.85334228442, 2191.85384798669, 
    2085.90431975464, 1697.12502302956, 1382.71016910742, 1348.56803552316, 
    860.452486946417, 643.441300007261, 2575, 2575, 2733.6222650195, 
    2733.6222650195, 2412.05612356136, 1938.91525080162, 425.785466617812, 
    100, 50, 40, -0, -0, -0, -0, 70, 90, 90, 90, 60, 60, 50, 50, 50, 40, -0, 
    -0, 40, 40, 40, 40, 40, 40, 40, 40, 50, 50, 50, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 160, 200, 210, 210, 210, 210, 180, 180, 180, 180, 120, 130, 
    130, 273.571165179653, 403.762466065914, 403.762466065914, 
    300.795080765481, 253.361404418945, -0, -0, -0, -0, -0, -0, -0, 2650, 
    3136.21196916827, 3587.10089597892, 3568.02712161929, 3485.03924236103, 
    3570.968181961, 3570.968181961, 3475, 3475, 3770.27681549167, 
    3804.20884127836, 3818.34664805503, 3833.86320691084, 3838.63240500181, 
    3831.86611713263, 3819.94639838263, 3820.04504627689, 3794.47607643191, 
    3761.37219263387, 3724.08007960673, 3701.89559479963, 3597.45201958195, 
    3258.47289616752, 2699.64487971633, 910.811933622343, 564.730534766639, 
    90, 120, 120, 120, 100, 90, 80, 70, 60, 50, 50, -0, -0, 60, 120, 120, 40, 
    100, 403.464575946532, 2775.47228438504, 4299.28965472685, 
    4299.28965472685, 4197.21482130183, 4041.92117523405, 3315.56322004115, 
    3722.71950624807, 3827.34670993386, 3778.44972539104, 3370.47502403535, 
    3599.39460145397, 3559.69632748161, 3330.36483743064, 3152.44393187334, 
    2598.56206036633, 2132.86569646581, 240.561416625977, 220, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 0, 50, 50, 90, 110, 110, 100, 100, 100, 50, 50, 
    50, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 130, 
    180, 354.314711364142, 1571.64007188392, 2533.60521475895, 
    2898.267022384, 3151.75548001105, 3357.94205220708, 3549.16147210279, 
    3588.58644662894, 3621.67621567091, 3701.9733920471, 3659.7172737033, 
    3582.49631833286, 3182.47995995106, 3355.18409166942, 3355.18409166942, 
    3350.64282558898, 3319.04233238735, 3301.59879305118, 3114.0753941246, 
    3036.92803911732, 2931.55586346119, 2611.08858516269, 2351.73791517767, 
    2250, 2250, 2250, 2250, 1575, 1575, 2922.03245664585, 2796.370519465, 
    2734.18647229723, 2872.01085829926, 3049.20974723112, 2836.44961797368, 
    2892.75569906168, 2198.9992449361, 1752.48889073994, 1422.89298557231, 
    1382.71016910742, 1327.67149942982, 953.492934812285, 583.651789906345, 
    375.311052633249, 334.226171713491, 1958.61565392935, 2412.05612356136, 
    2412.05612356136, 1938.91525080162, 1260, 140, 50, 40, -0, -0, -0, -0, 
    70, 90, 90, 90, 70, 130, 130, 100, 80, 60, 40, 40, -0, -0, -0, -0, -0, 
    -0, 40, 40, 60, 60, 60, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 150, 210, 210, 60, 60, 60, 80, 130, 130, 130, 130, 
    258.756995909204, 397.117183964076, 397.117183964076, 300.795080765481, 
    253.361404418945, 230, -0, -0, -0, -0, -0, -0, 2650, 3136.21196916827, 
    3568.02712161929, 3619.97389280298, 3485.03924236103, 3645.80682296714, 
    2442.6351058245, 1361.25975456197, 1579.67913375553, 3492.22280613679, 
    3701.68394692948, 3723.53886040094, 3773.69630568919, 3778.56284463689, 
    3814.13762999362, 3810.15910051528, 3811.08639295816, 3780.11789251868, 
    3740.72053597807, 3651.25015576531, 3274.45431670607, 2792.94869413153, 
    2630.27082205566, 180, 90, 90, 70, 90, 90, 80, 60, 60, 70, 70, 60, 50, 
    50, 70, 70, -0, -0, -0, -0, -0, -0, 100, 277.81534583022, 
    1754.4978841276, 3563.38255895111, 3563.38255895111, 3886.32976136971, 
    3886.32976136971, 3768.98779523247, 3783.16209905289, 3370.47502403535, 
    3370.47502403535, 3310.54322079629, 3261.20191465651, 2950.18284670323, 
    2309.17049991587, 643.556509060874, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 
    40, 60, 70, 80, 80, 90, 130, 140, 140, 130, 110, 80, 50, 50, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 180, 
    347.076139754556, 1998.58466378541, 2550.05190084888, 2859.94936230679, 
    3065.78548661781, 3286.00582782789, 3397.81617292101, 3488.66696834613, 
    3559.00624022418, 3608.98447769352, 3594.82977468166, 3452.52294044408, 
    3165.67357260236, 3112.63703106383, 3229.16288230858, 3350.64282558898, 
    3350.64282558898, 3359.05996309295, 3251.50170982941, 3238.18661629221, 
    3239.62530356273, 3122.78417752479, 3018.43148228355, 2555.69073555914, 
    2600.76983910411, 2345, 1975, 1975, 1975, 1975, 1425, 2507.5383483869, 
    2590.44345164368, 2734.82468817604, 2734.82468817604, 2836.44961797368, 
    3013.28614018553, 3033.85691278702, 2520.89403247056, 1863.26486472144, 
    985.734188349197, 955.428512809224, 1028.12928743958, 1028.12928743958, 
    990.145382927256, 270.610395222517, 150, 1673.18639959909, 
    1744.99605456957, 1744.99605456957, 1450, 1450, 40, -0, -0, -0, -0, -0, 
    70, 100, 100, 90, 80, 160, 160, 100, 80, 60, 40, 40, -0, -0, -0, -0, -0, 
    -0, 40, 40, 60, 90, 90, 40, -0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 40, 60, 60, 60, 60, 80, 130, 130, 130, 80, 190, 
    190, 170, 230, 240.561416625977, 240.561416625977, 120, 120, -0, -0, -0, 
    -0, 1350, 2844.6812571536, 3561.69907888819, 3561.69907888819, 
    3667.30509396827, 3490.35861655747, 2721.47223558249, 879.519343522738, 
    1684.04821561044, 3449.74919381534, 3470.10446188743, 3643.26774605444, 
    3643.26774605444, 3723.94568644628, 3728.98708133924, 3743.71183741367, 
    3721.27612304688, 3635.74941441696, 3284.82502657356, 2027.15106440345, 
    1421.65066047166, 370.154968261719, 370.154968261719, 130, 90, 90, 70, 
    70, 60, 50, 40, 40, 40, 40, 40, -0, 40, 70, 70, -0, -0, -0, -0, -0, -0, 
    100, 120, 140, 434.506022506018, 2332.75184361446, 3886.32976136971, 
    3886.32976136971, 3728.47671309042, 3549.7718750312, 3325.30062871749, 
    3325.30062871749, 2350.47681531575, 580.953491210938, 120, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 60, 80, 100, 100, 140, 150, 150, 130, 130, 140, 
    140, 130, 110, 80, 50, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 70, 170, 200, 1505.30024395573, 2425.71640768107, 
    2892.74505391147, 3100.32955893831, 3298.5618572555, 3287.80265268597, 
    3452.12812063305, 3458.3860302721, 3521.23157272932, 3536.10513914793, 
    3511.52402161935, 3476.87534425697, 3046.40560449008, 2738.15984583387, 
    2336.44039457858, 1864.18421823244, 2291.69187060417, 2670.99835930147, 
    3045.20248898006, 3128.15800038721, 3191.4755438382, 3195.90575871542, 
    3045.18973674089, 2980.66369488839, 2789.99582443548, 2606.89891429553, 
    2084.81303675708, 1975, 1975, 1975, 2169.02571952265, 1250, 1250, 
    2538.19604143944, 2722.6670877433, 2747.53212984665, 2900.2212400336, 
    2950.79436541311, 2919.8810768915, 2803.27663432128, 1717.69620672921, 
    738.966326273315, 1028.12928743958, 1065.54253797799, 1065.54253797799, 
    904.938022320088, 1186.84674527791, 1620.49673776301, 1768.2511908783, 
    1853.22008011058, 1450, 1450, 550, 550, 550, -0, -0, 60, 90, 130, 130, 
    120, 90, 190, 190, 50, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 
    60, 90, 90, 50, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 0, 240.561416625977, 240.561416625977, 230, 170, 100, 40, -0, -0, 60, 
    273.939235201579, 273.939235201579, 1053.17080285732, 2909.58635466928, 
    2951.71804149039, 2725.92853185723, 879.519343522738, 1684.04821561044, 
    3232.33867116081, 3323.75075739095, 3525.85775440526, 3643.03354628189, 
    3626.23218988866, 3601.16364921392, 3565.60136707275, 3226.57912363618, 
    3183.4956596064, 889.665641916594, 220, 140, 140, 110, 80, 70, 70, 60, 
    50, 50, 40, 40, 40, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 140, 140, 140, 120, 703.622538502745, 1213.73123434353, 
    1213.73123434353, 886.372088374374, 190, 150, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 60, 70, 100, 120, 140, 140, 150, 150, 150, 150, 150, 150, 150, 
    150, 150, 150, 70, -0, -0, -0, -0, -0, -0, -0, -0, 0, 120, 130, 130, -0, 
    -0, 60, 140, 180, 495.553629324057, 2039.13708314157, 2653.23052356179, 
    2907.115813202, 3065.78548661781, 3209.08194476896, 3287.80265268597, 
    3365.87836070389, 3430.78369401996, 3436.78816179894, 3425.97525623984, 
    3344.08171346483, 3230.93472926365, 3024.25397013054, 1942.85666763389, 
    782.38613351541, 765.980534677751, 750, 1356.0479406577, 
    2217.93267754086, 2699.35981519013, 2897.39251474069, 3038.49977064318, 
    3038.49977064318, 3046.67219463079, 2867.2758478028, 2703.0180673694, 
    2425, 2345, 2345, 1975, 1975, 1650, 1150, 985, 1050, 2431.55357345772, 
    2431.55357345772, 2595.56264574722, 2851.4588605582, 2790.42241257628, 
    2739.31048314251, 2565.82107686251, 1746.10063093739, 1245.93956499816, 
    1245.93956499816, 1163.82967487713, 1186.84674527791, 1368.44640917695, 
    1550, 1550, 1453.4565641416, 550, 1020, 1020, 775, 775, 775, 170, 90, 
    130, 130, 120, 110, 230, 230, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 90, 90, 50, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 230, 230, 230, 170, 100, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 987.570687765621, 1701.57221492236, 1740.00641417535, 
    2505.66105875573, 3093.22976460623, 3350.94250192195, 3139.62898537683, 
    2761.26582881083, 1526.82351844784, 964.799081546249, 210, 150, 130, 120, 
    90, 70, 40, 50, 50, 40, 40, 40, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 60, 70, 100, 130, 140, 140, 150, 150, 
    150, 150, 150, 150, 150, 150, 150, 150, 80, -0, -0, -0, -0, -0, -0, -0, 
    -0, 0, 120, 130, 170, 170, 200, 349.182690022309, 385.10121627728, 
    402.920754002841, 1126.63468249971, 2244.94241304162, 2598.30588722267, 
    2847.86352519875, 3012.44647037929, 3025.84194098294, 3108.5515180004, 
    3189.3087968145, 3259.13596493354, 3178.01283242697, 3065.78548661781, 
    2793.19719441086, 852.387088436488, 750, 120, -0, -0, -0, 
    552.840928865755, 1669.40156738965, 2148.26748651873, 2722.17761503025, 
    2937.59445353656, 2970.3620503418, 3014.56197902863, 2966.59084780835, 
    2425, 2425, 2345, 2345, 1975, 1975, 1650, 1350, 1350, 750, 750, 
    2036.36583307369, 2392.59583693207, 2587.48370053763, 2613.87977045527, 
    2549.01296136195, 2581.469500778, 2399.33186253102, 2399.33186253102, 
    2156.50980782973, 1840.89495099944, 1332.02543925047, 433.480353529111, 
    433.480353529111, 398.222505894324, 1020, 1020, 1020, 1020, 1020, 775, 
    775, 315, 0, 50, 130, 130, 110, 280, 280, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 0, 90, 90, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 170, 170, 90, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 70, 341.681821791071, 459.705153092628, 1131.9972401, 
    1131.9972401, 230, 190, 190, 160, 130, 120, 90, 70, 70, 50, 50, 50, 40, 
    40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 60, 70, 100, 130, 130, 140, 150, 150, 150, 150, 150, 150, 150, 
    100, 150, 150, 100, -0, -0, -0, -0, -0, 120, 120, 120, 120, 0, 130, 170, 
    170, 200, 349.182690022309, 385.10121627728, 460.538333080999, 
    1126.63468249971, 2193.13134777476, 2497.79652304161, 2692.17479494406, 
    2766.11152576309, 2795.31339759631, 2859.14438290328, 2965.24585782355, 
    3051.66037556653, 2885.38761804585, 1122.04064158262, 90, -0, -0, -0, -0, 
    -0, -0, -0, 550, 1920.91466207994, 2283.16401392661, 2492.94202824221, 
    2689.32411915296, 2842.4709468483, 2963.25480638061, 2345, 2345, 
    2345.48893969076, 2345.48893969076, 2126.69032951841, 1975, 1650, 1350, 
    1350, 850, 625, 1776.29559766656, 1812.3913446252, 1828.98287007791, 
    2142.94305978855, 2256.29431956149, 2319.9650789929, 2402.28382303851, 
    2399.33186253102, 2156.50980782973, 1840.89495099944, 1332.02543925047, 
    1150, 1150, 1150, 1150, 1150, 1020, 1020, 1020, 775, 775, 555, 
    557.934816991644, 200, 190, 210, 306.854010939725, 315, 315, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 90, 90, 90, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 100, 100, 90, 90, 90, 80, 50, 50, 40, 
    40, 40, 40, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 0, 70, 110, 140, 140, 130, 130, 130, 100, 40, 40, 
    100, 150, 150, 150, 150, 150, 150, 120, 120, 120, 120, 120, 120, -0, -0, 
    -0, 40, 40, 200, 274.560153501074, 460.538333080999, 1026.20860352967, 
    1421.0844711913, 1945.86711125925, 2380.214934007, 2453.65729009859, 
    2498.81165072749, 2527.807907711, 2540.47219367443, 2560.50379625668, 
    902.548483592609, 80, -0, -0, -0, -0, -0, -0, -0, -0, 110, 
    927.325982817347, 1796.45180622346, 2262.30219542944, 2274.12435092751, 
    2517.89385451306, 2734.33305998327, 2325, 2325, 2445, 2445, 
    2126.69032951841, 1975, 1669.7918181657, 1350, 985, 850, 550, 850, 
    1295.13488807675, 1339.65597605745, 1407.11310991943, 1606.89026335985, 
    1501.13942068031, 1841.30202097234, 2003.48836241176, 2056.95442663863, 
    1714.91765841599, 1209.74457092999, 1150, 1150, 1150, 1150, 1150, 0, 220, 
    475, 665, 665, 665, 1230.63414908473, 1230.63414908473, 864.651908564696, 
    640.635796632762, 474.92932486295, 315, 315, 80, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 90, 90, 90, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 70, 70, 80, 90, 90, 90, 80, 50, 50, -0, 
    -0, 40, 40, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 70, 70, 70, 70, 70, -0, 0, -0, 40, 40, 
    150, 150, 150, 150, 150, 150, 120, 120, 120, 120, -0, -0, -0, -0, -0, -0, 
    -0, 200, 255.152682383823, 270.610395222517, 456.840119440437, 
    862.448801342034, 1101.54602050781, 1627.20530666218, 1510.5853986913, 
    1409.84761277743, 1140.0801035984, 1140.0801035984, 230.074079547746, 70, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 90, 295.080183068428, 
    672.610825193284, 988.430036210461, 1937.91618805368, 2327.55673646024, 
    2325, 2325, 2445, 2445, 1975, 1971.1252066308, 1603.75281234831, 
    1365.7259344605, 985, 850, 850, 360, 360, 130, 70, -0, -0, 160, 
    315.148167399048, 662.955744949388, 1015.43771631363, 1015.43771631363, 
    473.476856554405, 378.652649329146, 446.606818287788, 450, 450, 450, 
    1643.4700950865, 2191.85384798669, 2522.44978660907, 2720.47512900157, 
    2702.31914186808, 2278.74635877007, 2089.38717901443, 1894.67591673689, 
    1532.96987738013, 1269.04766891606, 1269.04766891606, 1266.495546177, 
    642.352012364348, 230, 230, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    60, 60, 60, 60, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 70, 70, 70, 70, 80, 80, 40, -0, -0, -0, 
    -0, 40, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, -0, -0, -0, -0, 150, 
    150, 150, 100, -0, -0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 200, 
    311.603361361248, 310.52111384608, 353.773462632349, 359.117883173557, 
    721.308576036746, 736.670011762329, 736.670011762329, 736.670011762329, 
    304.134860603366, 140, 140, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 240.561416625977, 512.11091991334, 567.259843400989, 
    454.928195661354, 412.039822587801, 1497.18885950087, 1525, 1850, 1975, 
    1975, 1869.08706140525, 1550, 1050, 985, 985, 850, 360, 360, -0, -0, -0, 
    -0, -0, -0, -0, -0, 130, 220, 406.119789545056, 464.592428298097, 450, 
    450, 450, 2508.73874682691, 2784.05091232516, 3324.67999180097, 
    3125.43845649506, 3028.42611199966, 2847.22129266753, 2680.70765380889, 
    2597.31853312973, 2695.68937243938, 2106.93111379636, 1514.91714683636, 
    1266.495546177, 769.252552142694, 315.947316370387, 253.481433726992, 
    280.69671643634, 280.69671643634, 120, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 0, 60, 60, 60, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 
    -0, -0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -0, -0, 150, 150, 150, 150, 110, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 294.462890625, 345.517620388024, 
    425.785466617812, 650, 650, 650, 650, 650, 304.134860603366, 140, 140, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 260.314406253604, 
    326.990295410156, 391.452790222659, 412.039822587801, 627.95605812208, 
    985, 985, 985, 1050, 1150, 1150, 985, 985, 985, 985, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 130, 230, 444.398354275868, 839.197632807641, 
    803.625015916513, 990.840076931821, 1710.51683125018, 2508.73874682691, 
    2784.05091232516, 3227.30027818575, 3227.30027818575, 3221.27406198298, 
    3132.87602851633, 2989.36978048171, 2758.41088867188, 2515.78865629088, 
    2106.93111379636, 1514.91714683636, 1170.69263733482, 853.311387721143, 
    601.126073361421, 452.162459867855, 370.154968261719, 303.675919446708, 
    253.361404418945, 180, -0, -0, -0, -0, -0, -0, -0, -0, -0, 60, 60, 60, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 70, 70, 90, 90, 90, 90, 90, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 40, 
    40, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -0, -0, 150, 150, 150, 140, 110, 80, 70, 60, 50, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 312.079411495152, 345.517620388024, 
    468.074651616026, 650, 650, 650, 650, 382.223549174068, 294.462890625, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 985, 985, 985, 985, 985, 985, 1150, 1150, 985, 985, 985, 985, 
    985, 985, 985, 985, 785.185864282479, 253.361404418945, 305.503815291048, 
    326.990295410156, 370.154968261719, 773.951732148875, 1269.22395354106, 
    1402.35755290213, 1434.38824130697, 1558.49494612998, 1968.74497618778, 
    2706.27898331863, 3119.48440468526, 3240.7532773992, 3316.089559151, 
    3316.089559151, 3298.92759924097, 3088.07937618705, 2801.95133390926, 
    2344.17074520305, 1858.95236938763, 1561.48649587801, 1295.28082830596, 
    1027.18030769947, 814.848493014397, 659.102485947224, 527.263499343292, 
    425.785466617812, 344.34145084718, 258.574971126863, 190, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    70, 70, 90, 90, 90, 90, 90, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 60, 70, 70, 60, 50, 50, 50, 
    50, 50, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -0, 0, 150, 150, 140, 120, 100, 80, 70, 60, 50, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 360, 650, 650, 650, 650, 650, 
    347.659013195108, 270.610395222517, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 985, 985, 985, 985, 985, 
    1150, 1250, 1250, 1250, 1250, 1250, 1250, 1250, 1250, 1250, 
    785.185864282479, 811.773264009637, 850, 985, 1376.85269972816, 
    1535.46723323395, 1593.65386490985, 1680.8959319038, 1595.01098365763, 
    1742.72300524765, 2093.93249846243, 2695.6351373206, 3128.81661835894, 
    3330.82968769996, 3352.96750468838, 3352.96750468838, 3305.56315048051, 
    3134.26582347578, 2804.18770969183, 2324.6048995306, 1977.87843105849, 
    1765.08952739146, 1623.26682563758, 1478.68884277344, 1370.75672921834, 
    1261.50832329805, 1053.97168159182, 828.804923928544, 645.565741453072, 
    518.825939934596, 394.762851248428, 260.169551150474, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 90, 90, 90, 80, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 0, 70, 70, 70, 70, 70, 70, 70, 60, 60, 60, 
    50, 50, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -0, 0, 130, 130, 120, 110, 90, 80, 70, 60, 60, 60, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 360, 727.324662119998, 
    769.370730169722, 715.749076320971, 650, 650, 315.132705902373, 220, 150, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 985, 985, 985, 1150, 1250, 1250, 1250, 1250, 1250, 1250, 
    1350, 1350, 1350, 1350, 1186.76023600862, 850, 985, 1587.46305206827, 
    1653.69654712884, 1844.06477164239, 1851.13181259539, 1843.76282182733, 
    1896.23804707559, 2128.81879267655, 2616.32940893906, 3036.95865082194, 
    3243.30844403998, 3352.96750468838, 3377.08684414702, 3251.18141171095, 
    3019.87493996887, 2880.95234280607, 2743.84269999944, 2585.48344395201, 
    2447.70420703037, 2373.21388589408, 2312.62795999355, 2225.91588172602, 
    2140.71961250211, 1988.95597976277, 1720.9273974684, 1377.04333299493, 
    1090.21136179539, 834.852193654603, 668.612315318128, 548.869147973844, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 90, 90, 90, 80, -0, 70, 70, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 0, 0, -0, -0, -0, -0, -0, -0, 50, 50, 40, -0, -0, -0, -0, 
    -0, -0, -0, 90, 90, 90, 80, 80, 80, 80, 70, 70, 70, 70, 60, 60, 60, 50, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -0, -0, 110, 110, 110, 100, 80, 70, 70, 60, 60, 60, 60, 50, -0, 
    -0, -0, -0, -0, -0, -0, -0, 803.625015916513, 929.111551662542, 
    1030.74435225841, 988.794565216995, 785.824844346955, 650, 
    443.291929206742, 326.990295410156, 230, 180, 150, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    985, 1150, 1150, 1250, 1250, 1250, 1250, 1250, 1350, 1350, 1350, 1350, 
    1197.85510992233, 850, 985, 1548.34750358411, 1653.69654712884, 
    1749.05741301969, 1847.82542692495, 1843.76282182733, 1698.09865901325, 
    2045.7673284594, 2468.87289267096, 2758.41088867188, 2945.10028878918, 
    3074.75019739177, 3144.03443436363, 3113.14026990598, 3019.87493996887, 
    3023.83579722705, 3052.5961323357, 3052.5961323357, 3034.60478041413, 
    3009.76191201818, 2985.85331077544, 2928.23369421262, 2829.6937122446, 
    2709.91552700777, 2538.69138288981, 2352.43384710046, 2112.22198888281, 
    1806.79043396497, 1466.8320006904, 1154.89089676549, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 150, 150, 130, 100, 80, -0, 70, 70, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 40, 40, 40, 40, 40, 40, 40, 40, 50, 50, 50, 50, 50, 60, 
    60, 60, 60, 60, 90, 90, 90, 80, 80, 80, 80, 70, 70, 60, 60, 60, 50, 50, 
    50, 50, 50, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -0, -0, -0, 100, 100, 100, 80, 70, 70, 60, 60, 60, 60, 50, 
    -0, -0, -0, -0, -0, -0, -0, 826.40294604138, 1037.6739607335, 
    1207.58366640399, 1242.18725574051, 1242.18725574051, 924.771879268923, 
    707.724401746052, 521.503970643572, 370.154968261719, 253.361404418945, 
    200, 150, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 985, 985, 1350, 1350, 
    1350, 1350, 1350, 850, 850, 850, 1445.092417433, 1406.9586893066, 
    1360.51647313081, 1122.47006429062, 1150.36793302611, 1663.22082918686, 
    2081.45575837839, 2285.63699728708, 2451.64242545627, 2634.27398639561, 
    2787.93067079088, 2892.29798913686, 2956.46732737266, 3023.83579722705, 
    3052.5961323357, 3052.5961323357, 3034.60478041413, 3009.76191201818, 
    2985.85331077544, 3028.85909929022, 2960.15869697192, 2709.91552700777, 
    2538.69138288981, 2388.02812178583, 2223.1186307421, 2027.81403401561, 
    1749.98373454655, 1438.82490451903, 1060.28424242214, 747.785757239556, 
    527.632392811813, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 170, 170, 160, 150, 130, 110, 70, 70, 70, 70, 70, 60, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 50, 50, 50, 60, 
    60, 60, 60, 60, 60, -0, -0, 60, 60, 60, 60, 60, 60, 60, 50, 50, 50, 50, 
    50, 50, 50, 50, 50, 50, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -0, -0, -0, -0, -0, 80, 80, 70, 60, -0, -0, 50, 50, 50, -0, -0, 
    -0, -0, -0, 500.564715101512, 707.135493412933, 914.530756875361, 
    1159.63777823071, 1350.8037501805, 1350.8037501805, 1280.12060546875, 
    1082.27163169556, 833.426671384375, 530.481305895842, 376.703656250559, 
    294.462890625, 240.561416625977, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 481.129335533822, 625, 1550, 1550, 1550, 1550, 
    1382.7343320689, 850, 1150, 1703.47708947242, 1762.748729134, 
    1892.16770976963, 1864.8718962485, 1904.6182785089, 1998.56759676466, 
    2134.20198461711, 2232.79685000528, 2309.41042515317, 2407.70341051346, 
    2508.28550166627, 2659.21955672081, 2758.41088867188, 2824.45822310952, 
    2886.3238909981, 2916.12041268401, 2910.40331078037, 2875.72244429062, 
    2813.46000770178, 2733.34320657797, 2630.41912807999, 2513.60152271454, 
    2388.02812178583, 2223.1186307421, 2027.81403401561, 1749.98373454655, 
    1438.82490451903, 1060.28424242214, 747.785757239556, 527.632392811813, 
    326.990295410156, 294.462890625, 230, -0, -0, -0, -0, -0, -0, -0, -0, 
    190, 190, 200, 200, 200, 200, 200, 190, 180, 170, 160, 150, 130, 110, 90, 
    80, 70, 70, 70, 60, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 40, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 50, 
    50, 50, 50, 50, 50, 60, 60, 70, 70, 70, 70, 70, 70, 70, 70, 60, 60, 60, 
    50, 50, 50, 50, 60, 90, 130, 170, 240.561416625977, 327.576495897512, 
    425.785466617812, 568.633286553254, 696.95917008951, 803.625015916513, 
    803.625015916513, 785.088842857223, 988.027284546975, 1101.54602050781, 
    1175.87686660011, 1139.81969884721, 982.38670835712, 899.924293078008, 
    921.118951439175, 921.118951439175, 841.989871245989, 683.282409667969, 
    464.479332459468, 458.990158218235, 326.990295410156, 253.361404418945, 
    150, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, 80, 80, 70, 60, 
    40, -0, 0, 0, -0, -0, -0, -0, -0, -0, 500.564715101512, 727.293633152432, 
    835.240727725369, 1201.91758675948, 1397.8934598563, 1423.29106558656, 
    1365.67100370249, 1082.27163169556, 854.452506248158, 657.400413598855, 
    495.553629324057, 353.295952114701, 257.115871695691, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 340.863271979081, 625, 1550, 1550, 
    1550, 1550, 1550, 1853.0276970212, 2025.66391009482, 2149.03644382194, 
    2286.36020388254, 2340.47186396736, 2550, 2504.39123098378, 
    2550.46746974493, 2578.90297030026, 2613.17827467493, 2624.87826926281, 
    2591.23148115757, 2568.71871657567, 2563.19494692011, 2571.183032664, 
    2592.74384206647, 2607.17079182339, 2616.07178255952, 2610.75348948864, 
    2579.54504537522, 2517.55598443909, 2424.21428983262, 2292.02156964947, 
    2116.64898589393, 1935.05359591651, 1681.32135373606, 1430.8907167082, 
    1169.7028143082, 884.845586271986, 671.000513304544, 506.360868931452, 
    399.025221929836, 326.990295410156, 299.356564797915, 298.164369989564, 
    282.851637617016, 270.610395222517, 256.382279538765, 253.361404418945, 
    230, 230, 270.610395222517, 270.610395222517, 253.361404418945, 
    240.561416625977, 230, 230, 210, 210, 200, 200, 200, 190, 160, 140, 120, 
    110, 90, 80, 80, -0, 60, 60, 60, 60, -0, 60, 60, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 50, 50, 50, 50, 50, 
    50, 60, 60, 70, 80, 90, 100, 110, 120, 120, 120, 120, 110, 110, 110, 100, 
    90, 90, 100, 120, 170, 253.361404418945, 345.587278006649, 
    472.684962752598, 555.731769971044, 767.292996735217, 1071.19928901711, 
    1304.80212648975, 1520.05784710108, 1707.17007116932, 1898.87398704019, 
    2088.80583365255, 2207.43070126792, 2258.12471847336, 2300.27090037979, 
    2351.1489177105, 2416.2312260581, 2276.56471277279, 2151.20462207765, 
    2018.97412313362, 1935.05359591651, 1882.25407177628, 1625.37942473559, 
    1407.72620820993, 1183.75716287069, 947.683490287223, 699.68142462384, 
    460.400388089777, 335.933426786282, 210, 130, 80, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, 
    -0, -0, -0, -0, 80, 80, 70, 50, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 670.234803437528, 974.846966926886, 1323.29280203111, 
    1512.10721553113, 1628.75024508851, 1534.08762726743, 1280.12060546875, 
    1022.70207383598, 750.202524722497, 531.814170299302, 425.785466617812, 
    342.150168195457, 200, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 625, 1250, 1350, 1550, 1800, 2275, 2275, 2400, 2400, 
    2699.71580078802, 2743.12230426952, 2550, 3010.43513563493, 
    3050.55187678697, 3050.55187678697, 3015.45489250532, 3003.54029517127, 
    3001.91652501173, 2961.83629495136, 2922.43091550669, 2871.46030483447, 
    2801.80380587205, 2719.20276916313, 2636.71896248266, 2572.23905018542, 
    2483.70448495418, 2388.1114830509, 2272.66850188925, 2118.02783034573, 
    1892.33088850737, 1652.20512176987, 1362.64488153037, 1073.72588411079, 
    825.302267262008, 625.595028985913, 495.553629324057, 411.047557891161, 
    371.051375849609, 358.413526303035, 349.341867203907, 337.095958183899, 
    326.990295410156, 307.92271079354, 295.650179857504, 294.462890625, 
    284.457927263821, 284.457927263821, 281.739430630411, 276.055242314827, 
    270.610395222517, 257.602338016811, 253.361404418945, 240.561416625977, 
    240.561416625977, 240.561416625977, 240.561416625977, 230, 210, 190, 150, 
    140, 130, 110, 110, 100, 100, 100, 90, 90, 90, 90, 80, 80, 80, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 50, 50, 50, 50, 60, 60, 60, 70, 70, 80, 80, 90, 
    110, 130, 150, 180, 200, 230, 253.361404418945, 270.610395222517, 
    275.440795402962, 273.396719811597, 270.610395222517, 253.361404418945, 
    230, 210, 200, 210, 230, 275.78999695242, 346.370576212017, 
    452.757561680087, 620.172644977992, 824.025948084747, 1183.57514103089, 
    1601.44267506427, 1880.46616954808, 2191.85384798669, 2525.58248030263, 
    2818.49413699476, 3073.59127032374, 3147.51516519391, 3197.64054574195, 
    3268.75613891082, 3321.85181744882, 3387.2978515625, 3443.04625955465, 
    3263.28314814258, 3198.31352098043, 3128.03226210371, 3066.7830718901, 
    2894.60812630314, 2671.8000855559, 2515.32484999281, 2325.46015856573, 
    2121.30236846159, 1770.36559107882, 1511.50993818715, 1201.96116158727, 
    813.753409089106, 595.695209069526, 425.785466617812, 270.610395222517, 
    170, 120, 110, 90, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, 70, 70, 70, 50, 40, 40, 
    -0, -0, -0, -0, -0, -0, -0, -0, 740.340355651077, 906.369663649558, 
    1257.76587828429, 1532.40761254257, 1797.50000192078, 1791.55100588587, 
    1702.22097965625, 1551.25905326954, 1305.37437334944, 921.7500930649, 
    687.572057761914, 504.232736127317, 354.077714651925, 278.955612060767, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 440, 550, 1350, 
    1550, 1800, 2275, 2275, 2400, 2400, 2550, 2550, 2550, 3010.43513563493, 
    3050.55187678697, 3181.2430120949, 3325.55573945925, 3357.12713439233, 
    3373.16237321919, 3323.77623783941, 3259.86109088571, 3035.60588207748, 
    3053.71397430965, 2936.12047843126, 2737.55300427771, 2682.71781553726, 
    2544.64049533223, 2402.6626357, 2330.30423666223, 2159.75301982196, 
    1892.33088850737, 1652.20512176987, 1371.30354542422, 1051.65287963182, 
    755.070804720562, 547.038222772397, 425.785466617812, 383.181947928378, 
    378.913823138088, 358.413526303035, 349.341867203907, 337.095958183899, 
    359.519645284917, 359.519645284917, 344.068855603802, 326.990295410156, 
    312.739604373501, 299.604505237334, 294.462890625, 274.294991374762, 
    270.610395222517, 257.510545008055, 253.917739561212, 256.021158940257, 
    270.610395222517, 270.610395222517, 272.516651280041, 270.610395222517, 
    270.610395222517, 230, 200, 170, 150, 130, 120, 120, 120, 110, 110, 110, 
    110, 110, 100, 100, 100, 100, 90, 90, 80, -0, -0, -0, -0, -0, -0, -0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 0, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 40, 
    40, 40, 40, 40, 50, 50, 50, 60, 70, 70, 80, 100, 110, 130, 150, 180, 220, 
    260.052091702686, 326.990295410156, 402.959288247047, 495.553629324057, 
    594.669623417776, 683.282409667969, 757.095393577142, 806.244287746833, 
    858.518957875852, 884.576964855993, 855.982227568175, 775.51775435712, 
    702.119543579924, 580.953491210938, 468.917995872751, 408.016769926497, 
    452.230351094657, 540.391429821438, 660.729759136644, 819.915668782893, 
    1032.57133923449, 1306.39149491177, 1488.66510669365, 1647.32082619715, 
    2067.77830433115, 2566.462561134, 3008.04300838879, 3320.66093834101, 
    3530.86929959633, 3632.47839096141, 3677.50442723503, 3688.13533681493, 
    3688.25912670471, 3672.9391158193, 3635.13595054287, 3602.00370353162, 
    3552.92204794535, 3508.51591818216, 3423.62484426863, 3330.55713527612, 
    3222.78628089981, 3100.19583603584, 2915.38741300864, 2722.97604648154, 
    2530.76897796715, 2267.38762996469, 1964.00974015563, 1677.8047363475, 
    1378.34798372025, 1031.41014859526, 706.453525001649, 479.565009284697, 
    276.670683690594, 210, 180, 160, 190, 190, 170, 170, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, 50, 
    50, 50, 40, 40, -0, -0, -0, -0, -0, -0, -0, 731.305284933378, 
    751.107848512868, 1191.1341334413, 1511.59453177716, 1800.65346500796, 
    1935.24214734596, 1966.40812442881, 1935.05359591651, 1781.39475870434, 
    1401.08258628362, 1071.29302122932, 759.476599161267, 567.420972084093, 
    444.28606208837, 335.032432383896, 240.561416625977, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, 440, 440, 200, 1350, 1800, 1800, 1800, 
    2400, 2400, 2550, 2550, 2550, 2831.56451965241, 3045.38435153882, 
    3181.2430120949, 3325.55573945925, 3370.40211053634, 3357.12713439233, 
    3242.58343315526, 3094.90979439501, 3035.60588207748, 2957.63477271638, 
    2855.98422174122, 2737.55300427771, 2624.81643895845, 2547.62549979702, 
    2402.6626357, 2258.5838264837, 2060.10041984302, 1801.18709988714, 
    1479.3457784348, 1137.67734904855, 803.706570133992, 544.395290980734, 
    355.322329099469, 240.561416625977, 220, 220, 256.575971174801, 
    297.369886141245, 334.550944660301, 359.519645284917, 359.519645284917, 
    353.690241411623, 344.087273127727, 312.739604373501, 299.604505237334, 
    294.462890625, 273.675901664085, 258.610811099455, 253.361404418945, 
    253.361404418945, 256.337494414593, 270.610395222517, 278.274837030415, 
    294.462890625, 294.462890625, 275.4294110341, 255.008635896418, 230, 200, 
    170, 150, 140, 140, 130, 120, 110, 110, 110, 110, 160, 160, 150, 130, 90, 
    90, 80, -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, 40, 40, 40, 40, 40, 40, 40, 
    40, 50, 50, 50, 60, 70, 80, 90, 100, 120, 150, 190, 220, 
    258.250919121466, 313.863087363006, 382.638914182183, 443.400214549625, 
    580.953491210938, 708.227916203094, 852.696942436896, 957.594569218859, 
    1060.77410772889, 1144.68823785145, 1241.15861392874, 1382.58591003068, 
    1537.10177369615, 1644.23019250324, 1677.34157441696, 1614.62819219911, 
    1492.58057226416, 1280.31026753399, 1030.59974326674, 871.703357944241, 
    814.975822913979, 867.063045237582, 1043.92687902137, 1246.6980970536, 
    1379.89025109924, 1534.0907198193, 1616.51339321313, 1834.79423055321, 
    2139.43094985553, 2606.241538912, 3039.5258909797, 3377.03283736992, 
    3558.45640933334, 3705.20118109631, 3742.3029317394, 3731.2490901943, 
    3721.27612304688, 3693.50041291158, 3667.28813709262, 3639.91594128567, 
    3600.08599450516, 3562.01637151497, 3505.95454065229, 3444.66767689127, 
    3349.07179639197, 3236.71186330107, 3104.14964036313, 2941.34741374824, 
    2761.16062019149, 2570.09288574673, 2368.69171078783, 2016.56732516449, 
    1707.11379025988, 1388.39412766157, 995.657921235488, 671.720170035856, 
    456.086416439271, 306.548798837747, 253.361404418945, 230, 230, 230, 220, 
    200, 200, 200, 200, 200, 200, 180, 60, 60, 60, 60, 60, 40, 40, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -0, -0, -0, -0, -0, -0, 40, 40, 40, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 745.999442666131, 1080.98280073238, 1394.31002298698, 
    1618.23358199288, 1907.21835905127, 2016.21308051897, 2070.93268206792, 
    1997.74571087973, 1778.4170561061, 1426.98082375675, 1070.42803053122, 
    823.491038706779, 634.196052049806, 483.507116028614, 466.128446089024, 
    356.648661226347, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 190, 230, 240.561416625977, 258.804983708166, 279.809753322114, 
    409.351053691258, 1550, 1550, 959.883819285805, 1307.99582063521, 
    1939.71996273596, 2356.31845204454, 2678.39481047211, 2855.33118012431, 
    2973.44352261833, 3020.4213631239, 3005.20118284031, 2924.3006424619, 
    2799.67246820635, 2676.17170266009, 2563.77403103775, 2440.25029454267, 
    2256.77782566072, 2072.81556524677, 1898.5733788687, 1566.50944161561, 
    1236.00777490861, 929.207575843469, 654.35882933906, 443.159090132128, 
    280.082101557061, 150, 130, 120, 130, 160, 190, 240.561416625977, 
    273.969130965713, 302.817851499688, 326.990295410156, 326.990295410156, 
    300.987513757726, 283.058595042827, 271.325534992868, 270.610395222517, 
    253.361404418945, 241.006340868939, 241.618022983765, 253.361404418945, 
    260.003678951704, 275.057628536358, 294.462890625, 305.203959784114, 
    294.462890625, 280.442753050114, 270.610395222517, 240.561416625977, 210, 
    190, 160, 140, 130, 120, -0, -0, -0, -0, 160, 160, 160, 150, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 50, 50, 50, 
    60, 60, 70, 70, 80, 100, 110, 140, 170, 210, 253.858198514427, 
    326.990295410156, 397.478526070719, 501.757061013825, 645.536980273459, 
    816.12411308915, 974.381770106939, 1112.36946408882, 1200.03519000687, 
    1241.27192340827, 1295.81637428398, 1362.39560559433, 1409.38386061798, 
    1455.17209642491, 1556.05536299193, 1716.00694486155, 1846.5109779912, 
    1887.74484187567, 1856.00008420441, 1498.8668353644, 1280.31026753399, 
    1074.53798126922, 1057.79654852348, 905.494931873658, 1024.6102136827, 
    1143.62208487163, 1311.61123158576, 1431.42708146392, 1534.0907198193, 
    1561.50788915378, 1734.16939886011, 2060.12427157581, 2624.3745828857, 
    3039.5258909797, 3317.89582396114, 3600.3560490031, 3706.74733179282, 
    3761.71622798138, 3745.66393770172, 3729.41268306411, 3709.3749349656, 
    3683.96914465449, 3660.76362909274, 3631.4123928465, 3602.56040149214, 
    3552.4243945809, 3493.48104552771, 3418.43474249322, 3314.40664383961, 
    3218.93047220227, 3103.00074132086, 2971.27363312216, 2737.29735997612, 
    2421.60590958811, 2070.90253320992, 1857.95488959166, 1388.39412766157, 
    1075.26056281236, 671.720170035856, 456.086416439271, 306.548798837747, 
    253.361404418945, 230, 230, 230, 220, 200, 200, 200, 200, 200, 200, 180, 
    60, 60, 60, 60, 60, 40, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, 50, 50, 50, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, 650.401928125498, 768.615700761791, 
    1080.98280073238, 1361.3160207614, 1618.23358199288, 1799.65682390566, 
    1961.21186118932, 2049.31904775025, 1946.32981917209, 1771.18876253099, 
    1426.98082375675, 1125.72473767424, 893.771863160755, 655.543903201535, 
    561.205075386202, 478.811652934877, 409.670893392252, 326.990295410156, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 190, 200, 
    240.561416625977, 258.804983708166, 258.804983708166, 260, 1150, 1150, 
    473.962267290798, 745.645374046791, 1052.98078591201, 1741.76819224695, 
    2253.21712859568, 2555.77858989739, 2758.41088867188, 2859.21682377734, 
    2870.66114071581, 2794.55938081572, 2638.28427084426, 2466.66776221529, 
    2281.38180480176, 2055.27385727284, 1813.9567593421, 1502.23667670938, 
    1143.61952600912, 880.389692596403, 665.748897258852, 462.544490272626, 
    160, 160, 160, 140, 120, 110, 110, 120, 160, 200, 240.561416625977, 
    270.610395222517, 281.488977722084, 278.753266544652, 270.610395222517, 
    242.296219272358, 230, 230, 220, 220, 220, 230, 253.361404418945, 
    270.610395222517, 281.029706115772, 294.592914539463, 302.925544603904, 
    280.442753050114, 274.09539924958, 240.561416625977, 230, 200, 170, 140, 
    130, -0, -0, -0, -0, 180, 180, 190, 190, 190, 190, 190, 180, -0, -0, -0, 
    -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 40, 40, 40, 40, 40, 40, 40, 40, 50, 50, 60, 60, 60, 80, 100, 100, 
    80, 80, 70, 60, 50, 50, 50, 50, 50, 50, 50, 50, 50, 60, 60, 60, 60, 70, 
    80, 80, 90, 110, 140, 190, 258.674094037408, 355.673305113743, 
    457.879806896903, 610.37271745213, 803.625015916513, 960.982072973377, 
    1162.09990494995, 1380.4303175386, 1535.87196501642, 1706.61015014358, 
    1794.82861693066, 1811.46355017002, 1769.22061440166, 1705.65751932871, 
    1638.52558269776, 1579.11962490681, 1552.26950548763, 1569.90765728531, 
    1659.63114875163, 1776.07828355854, 1853.96367237828, 1883.41106941435, 
    1847.75624651178, 1498.8668353644, 1199.41972121507, 1074.53798126922, 
    961.685943548537, 905.494931873658, 1002.64616170553, 1358.45105611444, 
    1330.36461506646, 1431.42708146392, 1552.96762074626, 1697.12502302956, 
    1847.09346434451, 1994.024628862, 2619.92778699476, 3088.9953084882, 
    3393.97081755814, 3643.54431118564, 3706.74733179282, 3745.73687110675, 
    3733.86799756744, 3721.27612304688, 3704.3599546598, 3687.48916652107, 
    3670.12209195246, 3650.86209780324, 3616.76138730043, 3574.80303186463, 
    3524.89434724922, 3455.97498624459, 3374.0740161914, 3274.92274287688, 
    3139.00686090113, 2954.19907875682, 2737.29735997612, 2421.60590958811, 
    2070.90253320992, 1748.70330678741, 1207.56503172688, 860.299138310105, 
    581.945402746805, 413.34605803706, 240.561416625977, 200, -0, -0, -0, -0, 
    -0, 200, 200, 200, 200, -0, -0, -0, -0, -0, -0, -0, 40, 40, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, -0, 50, 50, 50, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    650.401928125498, 760.104453803964, 1007.30593644149, 1169.25137492511, 
    1347.49274657059, 1536.61229230337, 1738.76159929435, 1770.10681891696, 
    1752.01257144514, 1704.70274994468, 1422.63218234224, 1145.60908851293, 
    784.532990321551, 655.543903201535, 561.205075386202, 478.811652934877, 
    409.670893392252, 326.990295410156, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 140, 180, 180, 170, 190, 260, 985, 985, 
    340.656426619743, 659.399954205667, 988.256543017789, 1565.94411887364, 
    2080.92215123947, 2357.98781868385, 2497.92019608656, 2570.48267284005, 
    2553.57902067776, 2411.36275676989, 2171.64969086253, 1961.90730559062, 
    1726.01352781303, 1286.51300422885, 544.064664471434, 550.555495085408, 
    550.555495085408, -0, -0, -0, -0, 100, 100, 100, 100, 110, 110, 140, 160, 
    190, 230, 230, 240.808757233729, 242.762540884557, 242.762540884557, 230, 
    220, 220, 220, 220, 220, 220, 253.361404418945, 270.610395222517, 
    275.496262668161, 277.308206406078, 274.742245296696, 270.610395222517, 
    253.361404418945, 240.561416625977, 230, 200, 170, 140, -0, -0, -0, -0, 
    190, 190, 180, 190, 190, 190, 190, 190, 180, 150, 130, 120, 110, 90, 80, 
    -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 40, 40, 40, 40, 40, 40, 50, 50, 90, 140, 170, 230, 
    372.615849729007, 464.133391298049, 469.391843452785, 586.418672934597, 
    599.194339755176, 599.194339755176, 546.24946252735, 538.423378948757, 
    538.423378948757, 517.701987508925, 435.052138149071, 430.722542855762, 
    427.946618959138, 374.616590558731, 278.954521827072, 230, 200, 160, 180, 
    180, 170, 170, 200, 240.561416625977, 298.330492519539, 395.815116812934, 
    586.655702693574, 742.251012761651, 953.756994666289, 1206.56229789111, 
    1485.49676734753, 1749.802895462, 1979.51406332191, 2191.85384798669, 
    2317.8789064191, 2403.93887312184, 2439.79201373581, 2436.05360381317, 
    2388.56627991024, 2212.77875450164, 2018.11185158458, 1856.15504801054, 
    1773.46763932466, 1724.2550284077, 1739.90034572825, 1834.17585321371, 
    1964.94070964248, 2119.0639227999, 2250.02886404495, 2347.98967140887, 
    2429.87770268857, 2244.96685068884, 1973.91854867124, 1760.35756417515, 
    1552.37825322661, 1523.6705729086, 1550.60244303312, 1733.55386374204, 
    2007.60570557154, 2094.19277280754, 2099.92746673336, 2129.29616492049, 
    2304.8375897378, 2696.07716678962, 3022.6940466291, 3337.20696306588, 
    3530.1614926173, 3642.94753865868, 3706.74733179282, 3710.32901870444, 
    3702.71685886615, 3693.56079176367, 3682.23988335261, 3668.73768406053, 
    3662.91257659056, 3645.6849287167, 3624.14836612012, 3575.48408150325, 
    3508.81265217848, 3429.239393936, 3309.1506054086, 3125.98770444589, 
    3048.65931414596, 2619.27806915451, 2288.0202790286, 1935.05359591651, 
    1489.12011984674, 1029.10454879607, 785.36212229261, 568.725638774767, 
    335.339791072069, 253.361404418945, 170, -0, -0, -0, -0, -0, -0, 140, 
    140, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, 50, 
    50, 50, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    648.743041364228, 768.352969585599, 867.589439442949, 954.471508395082, 
    1059.98765901727, 1176.86558939327, 1280.12060546875, 1344.84607161839, 
    1387.94833348344, 1286.38987738748, 1101.54602050781, 818.572308786793, 
    692.670126841476, 546.82814691999, 428.422486586402, 408.564732693211, 
    342.670489852974, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 120, 130, 130, 130, 260, 294.462890625, 294.462890625, 
    445.101131314634, 705.177895136627, 1194.52738861836, 1728.19664916042, 
    2146.74735102891, 2401.35713244257, 2436.08225877235, 2436.08225877235, 
    2261.53944215224, 1952.07173440945, 1641.8151174535, 1310.6281687748, 
    884.286936685701, 500.949810013138, 434.337692337371, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 110, 150, 170, 180, 190, 190, 200, 200, 190, 200, 210, 
    220, 220, 220, 230.370433362452, 240.561416625977, 243.052055511561, 
    257.96221490754, 253.361404418945, 270.610395222517, 270.610395222517, 
    253.361404418945, 253.361404418945, 230, 210, 200, 200, 180, 160, 130, 
    -0, -0, -0, 200, 200, 190, 170, 160, 150, 160, 160, 160, 160, 150, 130, 
    120, 110, 90, 80, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 40, 60, 80, 130, 243.036298871737, 
    312.12666185763, 549.335733671926, 894.425912188474, 1126.87585245484, 
    1356.19244351782, 1697.12502302956, 1892.84426249011, 1935.05359591651, 
    2021.11439747525, 2133.00979470294, 2133.00979470294, 2065.19040661141, 
    2161.96448746878, 2158.92584818464, 2144.07942932536, 1951.95771290868, 
    1774.91970627194, 1624.79413172121, 1384.77302004162, 1145.97742286877, 
    998.724521339288, 942.839303029559, 942.839303029559, 975.308090998165, 
    1032.02687719003, 1047.12833221015, 1162.39464701667, 1364.6147688472, 
    1590.28068560614, 1770.59366916825, 1968.61500381946, 2164.87593113784, 
    2338.8126676486, 2475.00476466683, 2573.06259814254, 2636.5977695733, 
    2666.85485716857, 2676.60904837296, 2671.26997867223, 2644.72870507346, 
    2564.42513050625, 2507.23573136214, 2356.65645226589, 2141.61394913948, 
    2015.44664325579, 1969.09800205206, 2028.06328494988, 2166.56356633915, 
    2333.49546736369, 2519.48859747662, 2708.76024062579, 2902.80371766202, 
    3040.30911420228, 3051.07628284193, 3011.08064823015, 2954.4441530297, 
    2889.17773569071, 2853.9762170528, 2957.23784144686, 3016.56663507304, 
    3065.78548661781, 3116.41675767933, 3216.67572429997, 3302.4466145583, 
    3319.35405424186, 3387.83584540807, 3466.52630042236, 3609.24492297148, 
    3613.31169074272, 3681.44648714886, 3708.32998812269, 3704.20688084071, 
    3693.02409161359, 3681.50018698576, 3670.43498752795, 3655.65336628474, 
    3643.88849285889, 3635.91701007405, 3598.94902814104, 3552.40544326874, 
    3502.16046123346, 3390.06480738213, 3247.71515802895, 3065.78548661781, 
    2734.68292552688, 2400.25228664848, 1970.50803108465, 1558.34332613353, 
    993.485486809732, 859.903689219269, 634.200527195066, 481.844955883398, 
    337.981524384589, 220, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 40, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, 50, 50, 50, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 608.464289577926, 
    666.958947579646, 740.599266702126, 786.004623876037, 803.625015916513, 
    825.652865020005, 864.296044734264, 865.460373402569, 835.476647566044, 
    790.673592970221, 684.226613697935, 593.295100981229, 230, 
    316.681838305175, 316.681838305175, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 120, 130, 260, 
    270.610395222517, 448.48022272002, 724.095257013021, 1122.59547134346, 
    1824.94640982077, 2357.47423359491, 2447.41617413945, 2146.74735102891, 
    2142.65708382792, 1843.36937054681, 1526.5367710328, 1236.87912357229, 
    999.074528242111, 767.794040951113, 556.700812310455, 400.920645725987, 
    0, 0, -0, -0, -0, -0, -0, -0, -0, 150, 160, 170, 190, 210, 210, 200, 190, 
    190, 190, 190, 200, 210, 220, 220, 240.561416625977, 240.561416625977, 
    243.052055511561, 253.361404418945, 253.90313632398, 253.361404418945, 
    253.361404418945, 240.561416625977, 230, 210, 180, 180, 180, 170, -0, -0, 
    -0, -0, 200, 200, 200, 170, 150, 150, 140, 130, 130, 130, 110, 110, 100, 
    100, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 70, 90, 150, 294.462890625, 390.705959539201, 
    692.215092317248, 1140.41211931415, 1494.59280479774, 1812.86140918161, 
    2240.46275375746, 2495.05515824854, 2642.71052640899, 2858.63399383389, 
    2967.94937753973, 3011.54031464699, 3118.54047390421, 3188.83006107592, 
    3226.45738175629, 3253.37958712953, 3278.89779013413, 3244.89631879708, 
    3071.55858839859, 2844.13448092834, 2557.02529422544, 2236.99449055002, 
    1891.79046486513, 1806.33081420787, 1785.81015262688, 1804.45241910015, 
    1935.05359591651, 2126.08527422602, 2259.8820556722, 2393.33328492259, 
    2491.15864971465, 2568.35421833835, 2638.04728808083, 2698.24060412205, 
    2742.40738101575, 2728.51006613145, 2742.65882977991, 2774.62010291297, 
    2768.05420089671, 2768.69215084914, 2744.57080555431, 2694.49711305823, 
    2657.30985847516, 2564.97174997399, 2466.66776221529, 2332.79006777105, 
    2273.28000996592, 2291.51018470977, 2386.40083684147, 2552.52904741475, 
    2758.41088867188, 2931.35060413763, 3067.3953823442, 3182.62284205568, 
    3231.58905075312, 3247.90337878768, 3261.91800528107, 3281.59022246216, 
    3306.71273291279, 3364.5998427573, 3442.08801088385, 3499.04492747824, 
    3564.86885391403, 3602.40431797825, 3662.67099221188, 3680.64136001203, 
    3698.21855715122, 3707.59315336392, 3703.75277231426, 3703.75277231426, 
    3695.58693721432, 3708.25884189538, 3696.44652265528, 3682.5804606173, 
    3670.90907104489, 3650.40608457602, 3629.06479723475, 3609.07539478067, 
    3582.75507068107, 3551.59040991482, 3505.04657317512, 3442.66135641267, 
    3339.1713403875, 3212.99784255351, 2976.02390452647, 2652.99767854502, 
    2313.06207493044, 1855.64287562673, 1335.76855819199, 1040.30204180147, 
    718.814059113923, 547.855815430606, 432.463489744813, 379.006230482577, 
    326.990295410156, 260, 260, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 40, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, 60, 60, 60, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 355, 590.146896578851, 
    611.103393569932, 611.103393569932, 587.194412972082, 570.680195859608, 
    560.239164063725, 563.254939813162, 542.678415647161, 535.524435416612, 
    513.057907870593, 482.815369733355, 445.658883624293, 357.380974392673, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, 260, 803.625015916513, 1280.12060546875, 
    2126.13541124119, 2582.36945095434, 2732.47357220282, 2732.47357220282, 
    2453.85241194872, 2086.38600858991, 1649.5833965312, 1330.05783278736, 
    1143.40855925144, 1060.05655290513, 1089.37650943718, 1210.62253148252, 
    1210.62253148252, 1184.62941366193, 1019.18423529287, 819.152764322842, 
    601.657455055109, 353.863420002297, 279.932708996257, 160, -0, -0, -0, 
    160, 180, 180, 190, 210, 210, 230, 230, 220, 210, 220, 230, 230, 
    240.561416625977, 253.361404418945, 257.328451455065, 253.373558037017, 
    254.271075471227, 253.361404418945, 255.998752087478, 253.361404418945, 
    253.361404418945, 240.561416625977, 220, 190, 170, 160, 150, 140, -0, -0, 
    -0, 170, 200, 200, 180, 150, 130, 120, 110, 100, 100, 100, 100, -0, -0, 
    -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, 120, 150, 253.361404418945, 353.460424200313, 
    583.719420413804, 1005.21729959101, 1341.89622510073, 1794.80573415561, 
    2260.54302964885, 2556.19183403506, 2813.22870859709, 3025.22468062417, 
    3145.95906276657, 3248.95726000926, 3348.62964120234, 3416.37617986389, 
    3500.45288177527, 3586.46922432027, 3658.61372631208, 3674.31658462104, 
    3643.48623374301, 3614.13658471382, 3476.14562183279, 3195.55057793511, 
    2927.62868935534, 2627.04283754135, 2104.75884494956, 2018.84299766168, 
    1976.08443003085, 2021.95698612187, 2149.05133856437, 2366.03439272046, 
    2393.33328492259, 2576.8973521104, 2634.01676036914, 2668.97410961746, 
    2692.29218148299, 2711.72851427024, 2728.51006613145, 2742.65882977991, 
    2758.41088867188, 2777.12819206942, 2787.94652929257, 2758.41088867188, 
    2742.887495342, 2678.80796460938, 2583.82866940983, 2493.19874955104, 
    2432.65357947851, 2418.4292587733, 2476.26684585534, 2602.36464160173, 
    2711.03542847627, 2955.20194353262, 3118.37475441729, 3264.77478050232, 
    3344.17173765633, 3466.23464499217, 3521.67409164797, 3571.52829322419, 
    3607.85348927076, 3641.90407971691, 3616.31958712978, 3604.28005389117, 
    3609.62634528164, 3630.7902998903, 3642.20621925303, 3664.73074244941, 
    3676.9518824539, 3693.38524163613, 3701.58283785721, 3706.0176091502, 
    3703.75277231426, 3695.58693721432, 3682.52702205492, 3668.63843011615, 
    3646.11826928627, 3621.91704355809, 3597.5355638558, 3574.97395642297, 
    3545.57699417808, 3516.67998697932, 3462.9087218037, 3392.50984771998, 
    3314.04891325866, 3148.5762415536, 2943.82995913104, 2642.68817194385, 
    2225.56153981355, 1888.48560961376, 1389.32177481526, 870.812566374433, 
    712.116385197378, 497.061902752116, 373.927411828252, 340.097813448767, 
    332.544445714908, 335.113810933706, 260, 260, 260, 260, 260, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, 
    60, 80, 100, 100, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 275, 
    353.914097834774, 481.290348020289, 427.992237664823, 460.767133233811, 
    442.974617787455, 428.855618108036, 400.079867188216, 382.595557146494, 
    372.254622839032, 377.180137497491, 391.821507809983, 391.821507809983, 
    390.831769741334, 402.625561688495, 370.154968261719, 60, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    294.462890625, 439.5323942087, 669.394417592757, 1120.70967644776, 
    1728.68781619692, 2438.09049938469, 2837.87586800207, 3145.78713450315, 
    3196.91960401336, 3229.63102652618, 3172.55232775316, 3070.67540473893, 
    2833.57935041749, 2467.63957205786, 2145.44486040543, 1861.32393795486, 
    1649.51798239621, 1579.12820473293, 1641.42696075487, 1894.84798252525, 
    2081.17934824847, 2127.91460083486, 2034.85453768804, 1840.87064874875, 
    1497.08919901873, 1178.36956448635, 942.839303029559, 640.993608797265, 
    484.802857806091, 326.990295410156, 270.610395222517, 190, 180, 190, 200, 
    210, 240.561416625977, 257.974544071564, 259.550269505052, 
    254.051930773186, 253.361404418945, 230.218381528752, 242.698090995699, 
    253.361404418945, 257.831575931789, 270.610395222517, 274.392943448764, 
    256.772184724311, 254.284376626699, 253.361404418945, 253.361404418945, 
    253.361404418945, 230, 190, 180, 150, 140, 120, 120, -0, -0, 190, 190, 
    180, 180, 160, 130, 120, 100, 90, 90, 90, 80, 70, -0, -0, -0, -0, -0, -0, 
    -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 60, 90, 120, 150, 253.361404418945, 353.460424200313, 
    640.667022655988, 1005.21729959101, 1341.89622510073, 1898.93936000006, 
    2340.53855703729, 2720.47139960721, 3072.1897098128, 3205.11050159365, 
    3305.13020887407, 3391.6030590539, 3455.15482064659, 3526.60604088675, 
    3585.26840466372, 3690.53804268632, 3694.66573548973, 3825.49641880591, 
    3878.3827491877, 3898.19927275292, 3911.46592199956, 3929.56775979675, 
    3825.37804968986, 3662.77848394735, 3412.55468694531, 3266.68708095461, 
    2735.79022298594, 2406.44566185841, 2180.91487543271, 2113.38378623851, 
    2167.16449265821, 2240.39178075207, 2320.09198604235, 2395.22535868239, 
    2453.31048744988, 2487.71696924494, 2580.96375344861, 2747.67860919103, 
    2882.31445658508, 3002.1633395894, 3050.6609428487, 3050.6609428487, 
    3033.98257317619, 2943.81635169828, 2721.62087847678, 2629.50698206976, 
    2432.65357947851, 2418.4292587733, 2499.79288401649, 2579.80594220194, 
    2711.03542847627, 2886.88619229471, 3065.78548661781, 3232.94592927197, 
    3344.17173765633, 3411.17857447429, 3459.07718875999, 3505.56691751079, 
    3621.76148495931, 3534.28095912745, 3439.84700806482, 3370.17452723646, 
    3254.90115915924, 3312.90764873804, 3330.0345294349, 3401.94941159413, 
    3480.80878764717, 3540.70418600937, 3595.9379058951, 3650.09812693223, 
    3677.93638426655, 3686.24621020556, 3686.14776450835, 3662.161898645, 
    3635.89750576202, 3604.5273553541, 3557.76290145353, 3526.56197523079, 
    3462.32175857801, 3396.74971362457, 3327.54625254212, 3189.56284076819, 
    3039.48612645172, 2795.76972564816, 2466.66776221529, 2121.40608105452, 
    1582.67674183169, 1172.5267281532, 893.564255188506, 526.038319171484, 
    414.983853245102, 253.361404418945, -0, -0, -0, 243.308454873272, 260, 
    260, 260, 260, 260, 260, 260, 260, 260, 170, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 40, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, 80, 130, 140, 140, -0, -0, -0, 
    -0, -0, -0, -0, 274.845117211243, 274.845117211243, 275, 
    353.914097834774, 354.234202510594, -0, -0, -0, -0, 270.610395222517, 
    270.610395222517, 260, 256.568837991461, 308.080185882499, 
    315.168894565152, 370.154968261719, 370.154968261719, 375.615043814203, 
    60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    818.877302289799, 1087.75970114859, 1509.53200333237, 1858.28747552458, 
    2440.25999723938, 2800.7748310559, 3081.52808621816, 3512.53220339103, 
    3519.42896970071, 3106.06804381339, 3196.91960401336, 3211.6603987908, 
    3222.7295976185, 3369.12241375462, 3466.75243219316, 3490.84676590265, 
    3426.94810956923, 3313.96303253713, 3199.63179812877, 3038.69070866743, 
    2960.85587386228, 3095.50977563883, 3285.95095103942, 3506.33295873311, 
    3681.22581225308, 3410.24780968034, 3229.12156727096, 2991.73860753873, 
    2771.40808817195, 2089.55660761324, 1614.95944103935, 1073.81535447518, 
    686.426677985635, 507.924832834656, 377.963777043142, 280.443255069357, 
    272.550348900064, 277.020827026395, 240.561416625977, 257.974544071564, 
    257.974544071564, 254.051930773186, 253.361404418945, 230.218381528752, 
    242.698090995699, 254.373339392233, 257.831575931789, 270.610395222517, 
    270.610395222517, 256.772184724311, 254.284376626699, 253.361404418945, 
    253.361404418945, 240.561416625977, 220, 190, 180, 160, 150, -0, -0, -0, 
    -0, 190, 190, 180, 150, 140, 120, 100, 80, 70, 70, 60, 60, -0, -0, -0, 
    -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 60, 
    70, 70, 80, 90, 90, 90, 90, 90, -0, 326.990295410156, 640.667022655988, 
    877.812220692322, 1341.73235468056, 1898.93936000006, 2340.53855703729, 
    2720.47139960721, 3164.79169067092, 3252.72688596519, 3368.09141522975, 
    3464.24338248773, 3525.58340383296, 3566.27400315359, 3644.76826779743, 
    3690.53804268632, 3694.66573548973, 3800.86722739696, 3861.97167001236, 
    3933.00433933083, 3999.07353723049, 4051.71008218467, 4090.20884964745, 
    4107.17242865377, 4075.69955925464, 3950.11877117888, 3792.90894622602, 
    3486.80218914733, 3096.09950992822, 2698.33561345744, 2358.17458696484, 
    1800.34631665478, 1923.76762208145, 1945.73902683889, 2027.21331653448, 
    2206.44834097887, 2505.61268208849, 2747.67860919103, 2882.31445658508, 
    3191.39997947298, 3246.23319683816, 3195.480275874, 3011.68420788934, 
    2958.96995457857, 2721.62087847678, 2442.3589936877, 2264.98656743417, 
    2145.76030299765, 2072.21913804208, 2086.18534854595, 2144.77181589431, 
    2191.85384798669, 2303.85147691194, 2401.21935236911, 2477.32397706433, 
    2600.11995854808, 2730.28363473972, 2823.62630756041, 2867.56819361934, 
    2896.48866708312, 2909.19304694552, 2880.57056167062, 2865.78374428258, 
    2885.10894501737, 2944.02252590547, 3075.77710911778, 3180.77621829541, 
    3327.05403724501, 3466.74164359279, 3552.53632457235, 3619.49577799756, 
    3637.14186127867, 3641.50335189371, 3613.54933863364, 3557.20618613519, 
    3509.35233064936, 3399.2712199282, 3304.81686394154, 3207.22874953398, 
    3118.54219442689, 3021.04104537514, 2866.17177655651, 2734.82077507125, 
    2415.29925377456, 1998.91275290516, 1633.85288312462, 1105.35001959329, 
    813.650473379844, 533.017517030415, 343.35944223995, 230, -0, 0, 0, -0, 
    -0, -0, -0, -0, 260, 260, 260, 260, 260, 260, 210, 180, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, 40, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, 130, 160, 180, 190, 
    190, 190, 190, 190, 190, 190, 281.837540882536, 281.22746911677, 275, 
    275, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 60, 60, 60, 60, 
    60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 170, 
    270.610395222517, 314.914240448569, 313.310271860009, 315.682985951006, 
    294.462890625, 294.462890625, 301.595578836499, 278.78536923144, 
    415.597755064152, 560.243759428911, 560.243759428911, 557.376738196627, 
    393.924442507384, 589.693839058697, 727.078828114783, 894.441200537819, 
    1147.92650096056, 1478.68884277344, 1858.28747552458, 2440.25999723938, 
    2800.7748310559, 3081.52808621816, 3658.41417210777, 3690.86230456788, 
    3662.09455116272, 3540.17054838059, 3387.2978515625, 3331.84923728253, 
    3368.21947826924, 3412.35026896895, 3489.31323303213, 3572.69909673481, 
    3665.25503649167, 3636.32332297613, 3831.80920443467, 3894.57855617197, 
    3962.29956284468, 4004.49580516727, 4016.48314420348, 3976.65535848707, 
    3909.45330215862, 3811.16117676721, 3605.46005246838, 3330.5187217139, 
    3012.53048646793, 2539.20006374314, 2027.58463360333, 1554.57301743489, 
    995.820472691718, 771.299453450189, 580.953491210938, 386.029666896287, 
    281.391211542623, 240.561416625977, 220, 200, -0, -0, 170, 190, 220, 
    230.555413559682, 230.555413559682, 230, 230, 230, 230, 240.561416625977, 
    240.561416625977, 240.561416625977, 240.561416625977, 210, 190, 170, 150, 
    -0, -0, -0, 180, 180, 170, 140, 120, 100, 70, 60, 50, 40, -0, -0, -0, -0, 
    -0, -0, -0, -0, 40, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 50, 60, 
    70, 70, 80, 90, 90, 90, -0, -0, -0, 0, 406.359925346723, 
    551.415242288792, 890.823120821558, 1313.1913133105, 1790.82114614882, 
    2218.76328351277, 2765.16767326591, 2991.22918750725, 3234.37802382856, 
    3373.44165758673, 3445.68366771813, 3513.83099951363, 3564.75912725961, 
    3577.57940252971, 3620.41211356566, 3697.21228142653, 3802.17161208536, 
    3810.84267791777, 3901.46029653244, 3983.91882810885, 4089.73746919612, 
    4161.0535455802, 4204.1757877174, 4196.24113124406, 4173.36562818469, 
    4118.4304225315, 4040.65724421965, 3884.68938054716, 3615.10267109383, 
    3222.06164296295, 2779.08603219013, 2220.82201499243, 1821.84291160773, 
    1666.10264212361, 1833.56623108266, 2254.83727463316, 2766.24354816516, 
    3248.51956302137, 3339.56833750513, 3106.78148197433, 2798.91228302458, 
    2786.31229860041, 2688.86126610925, 2587.49528329936, 2469.06149207939, 
    2321.31551368568, 2146.09860875225, 2016.34327137457, 1953.97940182308, 
    1978.75156259833, 2039.4273001576, 2080.49612408751, 2117.96786231352, 
    2171.28843122793, 2218.5303227265, 2301.43940669891, 2376.33633610394, 
    2466.66776221529, 2478.06512421544, 2572.11829921267, 2685.96418407735, 
    2795.00547531013, 2940.54683180418, 3095.47235066755, 3252.02910491426, 
    3374.97899496882, 3479.6370825705, 3512.33786442701, 3538.64391563364, 
    3535.78525511552, 3521.17080275392, 3493.02628925964, 3425.31435417925, 
    3359.94086961717, 3215.80255471093, 3078.03910552024, 2976.83055312846, 
    2818.73340868766, 2671.59350367553, 2502.45723534672, 2431.20109108229, 
    2000.9756414966, 1726.87569316234, 1313.29207381333, 819.206390430797, 
    637.307466009187, 391.440737024218, 275.449219525778, 0, 0, 150, 150, 
    140, 140, -0, -0, -0, -0, -0, 253.361404418945, 260.232885305827, 
    279.941047508635, 270.610395222517, 210, 210, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 40, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, 160, 180, 190, 190, 190, 
    190, 190, 190, 190, 190, 190, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 60, 60, 60, 60, 
    60, 60, 60, 60, 60, 60, 60, 170, 270.610395222517, 315.144722500371, 
    350.109647966291, 524.393175092674, 670.452695519308, 651.045626288304, 
    1019.56582547217, 1412.36540794545, 1495.68533248076, 1673.10585149614, 
    2027.80399852673, 2124.85368531815, 2138.46186618661, 2016.86195561456, 
    1814.6668738844, 1832.12276656212, 2012.8670383515, 2218.45947187743, 
    2359.9075451784, 2466.66776221529, 2540.48050675678, 2627.27446009847, 
    3439.08217611943, 3892.62483912712, 3957.37137004362, 4005.07192445458, 
    3930.78377948827, 3829.10975550528, 3721.81113349996, 3636.22721715703, 
    3588.99669263828, 3550.89163849949, 3559.47192622344, 3636.32332297613, 
    3721.27612304688, 3815.09898822401, 3892.1651240078, 3913.80040559235, 
    3934.2093897203, 3944.74208646063, 3943.16116526523, 3887.36258704359, 
    3811.55621726925, 3746.04536021399, 3528.11067077002, 3280.8996256548, 
    2987.89760669541, 2448.10529720761, 1921.23361534842, 1280.27681411847, 
    902.448340886097, 528.578192805605, 307.63864562536, 254.830953535959, 
    230, 200, 0, 0, 150, 150, 0, 0, 190, 210, 210, 220, 240.561416625977, 
    256.052701911101, 270.610395222517, 281.916056595343, 270.610395222517, 
    240.652879150468, 240.561416625977, 210, 200, -0, -0, -0, 180, 180, 150, 
    130, 100, 70, 60, 40, 40, 40, -0, -0, -0, -0, -0, 40, 40, 40, 40, 40, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 40, 40, 40, 40, 50, 50, 50, 
    60, 60, 70, 70, 70, -0, -0, -0, -0, -0, -0, 271.645401849563, 
    409.132135696785, 719.474069671483, 868.33178372195, 1546.73315949337, 
    2006.310031948, 2466.66776221529, 2843.87184083013, 3154.16094269167, 
    3319.13462561449, 3441.53268582955, 3483.34663856035, 3531.14682435354, 
    3549.77844414838, 3564.88962295236, 3589.03700506861, 3707.83192654735, 
    3886.56279543994, 3913.62401631884, 4016.85964259101, 4111.33675788722, 
    4164.39289975305, 4218.30658323912, 4224.62108530328, 4218.80515262627, 
    4200.63707854396, 4173.06071698592, 4065.89147763595, 3805.62148167833, 
    3363.53270338954, 2929.55694961715, 2090.01804097267, 1586.09082961729, 
    1446.34171649125, 1697.12502302956, 2347.40439156871, 3202.10985206597, 
    3640.4053194002, 3776.60607965536, 3759.72537683854, 3701.60229704952, 
    3682.85805201113, 3654.81504552083, 3608.88801205444, 3538.42262733026, 
    3319.87922687201, 3187.54306736163, 3081.33642376911, 2969.26769216137, 
    2758.41088867188, 2490.63995477148, 2403.71881461167, 2160.3651235736, 
    2160.3651235736, 2118.10264843481, 2098.88851354745, 2150.84465657364, 
    2253.50773291903, 2373.53488390358, 2586.90962605929, 2780.22660113162, 
    2975.07734216279, 3148.88008976818, 3244.0588854032, 3294.94499601188, 
    3358.40021294387, 3321.78873854011, 3277.92802840983, 3297.58617806124, 
    3265.0656808654, 3226.12717003938, 3163.09371952099, 3101.802034057, 
    2983.19136915474, 2871.30927216656, 2675.82478066874, 2484.85453266054, 
    2207.28277645791, 1924.17207563043, 1660.58062581827, 1374.20120464878, 
    1106.68709340622, 803.625015916513, 599.085045466468, 411.081030778115, 
    294.462890625, 210, 180, 170, 190, 240.561416625977, 240.561416625977, 
    230, 210, 0, 0, -0, -0, -0, 259.147622653471, 270.610395222517, 
    281.539288532534, 243.250938789507, 210, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, 40, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, 150, 150, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 276.217709570817, 353.220940440763, 513.396551434776, 
    657.585517752349, 844.068959826272, 912.43346307374, 912.43346307374, 
    912.43346307374, 1019.56582547217, 1354.60121838794, 1495.68533248076, 
    1673.10585149614, 2062.2726048351, 2124.85368531815, 2124.85368531815, 
    2016.86195561456, 2327.35674966298, 3207.46954716297, 3389.67611398536, 
    3681.67676921833, 3851.31341095936, 3998.6508255509, 4094.32616517388, 
    4138.48238447995, 4160.07475422953, 4185.66304335665, 4190.38003822379, 
    4173.69117764016, 4141.71375740089, 4076.43135986316, 3963.97725785946, 
    3798.66020352789, 3601.88694739097, 3464.05182030659, 3531.37212857712, 
    3467.55845023642, 3505.55076251379, 3567.89424203948, 3652.57174219262, 
    3782.74920164584, 3835.61129240174, 3856.89416679282, 3882.70330666617, 
    3872.33528288144, 3858.46967937641, 3827.40332232789, 3800.41894892039, 
    3657.03545311729, 3508.36005183595, 3142.62519810312, 2618.51117059647, 
    2065.86463849345, 1459.39926458817, 881.746769308616, 547.928634565497, 
    391.819554384751, 230, 190, 140, 140, 140, 140, -0, -0, 210, 
    240.561416625977, 254.690634677367, 277.216246080049, 308.528093732103, 
    326.990295410156, 335.160141818363, 341.741732792962, 331.163117354916, 
    326.990295410156, 304.767920880624, 294.462890625, 240.561416625977, 230, 
    190, 180, 160, 160, 130, 100, 80, 60, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 50, 50, 60, 60, 70, 
    80, 90, 100, 110, 110, 100, 0, -0, -0, -0, -0, -0, -0, 612.993426996865, 
    1021.3680065325, 1567.98702210212, 2119.96910341317, 2516.13397592101, 
    2971.21221151367, 3165.00595924749, 3331.84341489287, 3439.14293422414, 
    3505.19762301191, 3555.14036966554, 3604.20075615975, 3638.75302742858, 
    3707.83192654735, 3835.40341406473, 3864.03557952878, 3947.10675653365, 
    4014.62566194123, 4143.31602868684, 4222.49619538953, 4244.48874936052, 
    4250.44706148513, 4247.12852941086, 4235.31711286058, 4213.2669670846, 
    4137.89289902809, 3830.62268473855, 3354.1879280524, 2705.55791144583, 
    2124.28280930517, 1851.47567699334, 1851.47567699334, 2347.40439156871, 
    3330.77064574532, 3640.4053194002, 3845.34456255063, 3840.60989617221, 
    3701.60229704952, 3682.85805201113, 3654.81504552083, 3621.03942530417, 
    3513.0040323912, 3319.87922687201, 3187.54306736163, 3273.78525989521, 
    2969.26769216137, 2905.47473234269, 2681.91370427122, 2385.52822665096, 
    2145.15087717583, 1990.31877981169, 1863.89483709364, 1786.80553725848, 
    1845.50686474166, 2001.8555956327, 2077.4953267121, 2321.18413157715, 
    2467.43830980293, 2629.90690013984, 2818.78293593666, 2874.80702311296, 
    2962.20018988894, 3032.58391235787, 3076.93083087286, 3142.04682900544, 
    3120.19277159522, 3151.49989745682, 3065.78548661781, 2965.94748047182, 
    2847.56423270318, 2715.76575906729, 2466.66776221529, 2252.17723327233, 
    1914.37341002397, 1597.73681867768, 1292.10481582081, 1005.78887797578, 
    812.240182820934, 652.055185909333, 532.495961873339, 427.27888805378, 
    370.154968261719, 210, 240.561416625977, 240.561416625977, 
    253.361404418945, 253.361404418945, 240.561416625977, 240.561416625977, 
    230, 210, 0, 0, -0, -0, -0, 210, 256.266061203684, 253.361404418945, 
    243.250938789507, -0, -0, 160, 160, 140, 140, 130, 120, 90, 40, 40, 40, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 60, 60, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 60, 60, 
    60, 60, 60, 60, 60, -0, -0, -0, -0, 160, 160, 160, 160, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    253.694527001745, 451.565025334818, 523.336000457975, 639.375049824849, 
    832.088692728572, 919.728072957004, 984.822755601026, 1078.83538088292, 
    1032.53495827018, 990.926651552624, 912.43346307374, 912.43346307374, 
    860.05589341834, 878.941961943347, 883.142757273458, 883.142757273458, 
    1037.81490360744, 1088.62728481282, 1230.58644327839, 1842.32822016647, 
    2327.35674966298, 3065.78548661781, 3401.32805302732, 3655.46631133256, 
    3877.883296679, 4013.09882186733, 4133.55510745616, 4202.74983823221, 
    4143.63231645383, 4286.77692440186, 4264.15830882231, 4239.28826293418, 
    4247.26980132354, 4248.41400909934, 4216.85843985815, 4146.24123084066, 
    3913.37312499509, 3804.1508567804, 3601.97448261392, 3508.51482283386, 
    3527.6514563427, 3554.6153735187, 3621.16924686764, 3692.17351340217, 
    3787.53084615104, 3838.25034340679, 3829.6886597642, 3824.68155239391, 
    3809.69880437688, 3786.58550845751, 3766.72252726767, 3657.03545311729, 
    3672.31929346352, 3466.00612885375, 3244.97996162897, 2886.70115750579, 
    2343.60389977792, 1843.38274278812, 1432.1212602246, 877.642270610953, 
    740.070188532561, 530.829233148352, 394.687149720632, 376.014418103491, 
    338.769934875539, 354.914484991669, 370.154968261719, 382.494920517763, 
    402.107685511792, 412.958443777673, 388.594568434013, 370.154968261719, 
    370.154968261719, 349.251617354072, 349.251617354072, 335.160141818363, 
    331.163117354916, 326.990295410156, 304.767920880624, 302.927479278211, 
    240.561416625977, 230, 190, 180, 150, 130, 100, 80, 60, 50, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 40, 40, 40, 40, 40, 40, 40, 50, 50, 50, 60, 60, 70, 80, 
    90, 100, 100, 110, 110, 120, 130, 150, 170, 200, 220, 220, 
    270.610395222517, 326.990295410156, 529.862069377942, 822.950314068296, 
    1243.53405244182, 1754.53313198731, 2355.97831102532, 2672.63025843132, 
    3097.61988263986, 3258.11731634505, 3455.13839148849, 3505.38071814127, 
    3575.93282055024, 3594.73924084198, 3620.90153331393, 3643.29464275893, 
    3677.68745337874, 3721.27612304688, 3799.76121975822, 3817.96801040771, 
    3985.41706626637, 4136.29872774845, 4187.59366937519, 4255.89010678795, 
    4269.43475900936, 4270.66574183747, 4268.30580065881, 4236.45630558452, 
    4146.69545196829, 3926.93128020243, 3436.77048822479, 2934.41232263827, 
    2414.63536381649, 1881.27957175938, 1809.3467990769, 2268.37418985841, 
    2711.67221115286, 2996.54212724084, 3128.87827662759, 3548.51460315015, 
    3680.00482152513, 3620.42457010305, 3426.46552363583, 3231.9092040979, 
    3159.40215489394, 3139.65929930514, 3079.98645637758, 2888.50964216107, 
    2733.98849245241, 2513.2647442035, 2272.71081886898, 2081.15193692109, 
    1960.38699829604, 1829.9749961303, 1824.69373663745, 1655.67673459809, 
    1495.14681483419, 1591.41939567992, 1655.4191074487, 1697.12502302956, 
    1884.82638787985, 1936.05277890654, 2148.41834656022, 2283.36071549481, 
    2466.66776221529, 2660.89113006489, 2741.35233309484, 2822.39902910171, 
    2854.86029206242, 2863.02044251099, 2714.92694543742, 2583.99144572579, 
    2299.19096021661, 2033.67187887465, 1665.15646602774, 1338.27048848948, 
    1022.23173134002, 812.468135231354, 645.566928438421, 528.707161081315, 
    459.555813956481, 408.863115322134, 376.61968325472, 359.212210479001, 
    210, 240.561416625977, 240.561416625977, 253.361404418945, 
    253.712853952849, 210, 210, 210, 170, 0, 0, -0, 80, 110, 160, 190, 200, 
    200, 160, 160, 160, 160, 140, 140, 130, 120, 100, 80, 40, 40, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 60, 80, 90, 90, -0, -0, -0, -0, -0, -0, -0, 110, 120, 120, 60, 60, 60, 
    60, 60, -0, -0, -0, -0, 160, 160, 160, 160, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, 0, 0, 0, 240.561416625977, 278.805401622913, 384.92780145636, 
    495.553629324057, 685.728964580604, 762.551465960489, 1013.82501230238, 
    1269.2904831834, 1349.11222683155, 1530.89956841899, 1602.36321850324, 
    1697.12502302956, 1702.70654183705, 1787.28703283309, 1800.26586416545, 
    1850.81574953952, 1906.96786125279, 1958.10839168436, 2080.88257438359, 
    2110.31079064119, 2222.13702751134, 2246.25488742347, 2216.45799940563, 
    2231.90170784877, 1890.01434411346, 1615.45454228832, 1418.36319946739, 
    1684.65545763003, 2108.88803690757, 2797.09038432379, 3329.30626315952, 
    3749.25325252889, 4016.92946026956, 4182.66226053133, 4254.27765638444, 
    4294.84358205526, 4272.81436378453, 4291.72756248286, 4274.95220244753, 
    4254.72849284889, 4245.18584436554, 4225.33653250624, 4156.8187125071, 
    4044.9471620807, 3844.850193842, 3732.08832513997, 3696.19307317385, 
    3479.99747543124, 3411.45455111962, 3411.22306593971, 3521.1424704068, 
    3562.00596585274, 3647.98037512899, 3690.5397705723, 3707.18594678493, 
    3700.59736967443, 3683.92963314129, 3620.08261066109, 3580.38280657087, 
    3450.00334072523, 3343.01470911514, 3112.84434017739, 2878.86324180866, 
    2510.0365471285, 2131.0501301521, 1728.86013420199, 1295.3402789618, 
    1034.11527402636, 813.912930067905, 644.772093499148, 536.125258972534, 
    354.914484991669, 370.154968261719, 382.494920517763, 393.356726825349, 
    393.356726825349, 388.594568434013, 370.154968261719, 370.154968261719, 
    349.251617354072, 350.724375667063, 333.282266163076, 330.643337493783, 
    306.973602951276, 300.839160325396, 260.007681549889, 240.561416625977, 
    200, 180, 140, 120, 90, 80, 60, 50, 40, 40, 40, 40, 40, 40, 40, 40, -0, 
    -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, 40, 40, 40, 40, 40, 40, 50, 50, 60, 70, 70, 80, 80, 90, 
    100, 100, 100, 110, 110, 120, 130, 150, 170, 200, 220, 253.361404418945, 
    296.331716767275, 396.259039671258, 570.088791309225, 722.526943397964, 
    1168.09269205588, 1519.14920238414, 2034.67733393124, 2466.66776221529, 
    2813.26470780158, 3076.93070443612, 3278.19747077479, 3402.47521936914, 
    3478.94771724321, 3530.22170256221, 3559.34898807307, 3604.69171201514, 
    3606.572411053, 3674.9512403301, 3729.08615771251, 3776.52727446498, 
    3811.50864663906, 3913.93678015072, 4065.89147763595, 4140.91597614515, 
    4246.4881370971, 4285.27927119633, 4291.01624335326, 4276.21627746928, 
    4275.43129579895, 4273.8930829705, 4258.43328291573, 4245.47746183157, 
    4224.49186497179, 4201.08781381872, 4145.9822750494, 4149.89924676527, 
    4170.67118068016, 4086.86252930586, 3669.6815452323, 3432.80491116969, 
    2964.38782913142, 2404.96579197073, 2495.922254205, 3081.75928412296, 
    3341.24045372438, 3235.72191068418, 3138.85465274671, 3065.78548661781, 
    2945.94105383276, 2690.03721974888, 2469.1876719985, 2267.93234548026, 
    2017.82638546261, 1907.72603424672, 1725.10420428374, 1616.19113114244, 
    1566.43825216009, 1504.10076503933, 1526.59731661951, 1506.09096290633, 
    1528.69450247657, 1556.78903584198, 1609.78670165883, 1733.72905239524, 
    1848.87321279065, 2027.8755404193, 2136.58170248376, 2233.5154994501, 
    2253.05991211617, 2080.92424694339, 1874.32821262216, 1645.6997278156, 
    1330.32728706004, 1131.53605951877, 879.231236315021, 741.165377978484, 
    559.55660092983, 495.553629324057, 412.199750718103, 379.252351912604, 
    370.154968261719, 336.903964974572, 326.990295410156, -0, -0, -0, -0, 
    220, 220, 220, 220, 230, -0, -0, -0, -0, 80, 110, 160, 160, 160, 160, 
    160, 160, 160, 160, -0, 120, 110, 110, 100, 80, 50, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 
    80, 90, 100, -0, -0, -0, -0, -0, -0, -0, 110, 120, 120, -0, -0, -0, -0, 
    -0, -0, -0, 180, 180, 180, 180, 180, -0, -0, 0, 0, 0, 274.827602371158, 
    253.361404418945, 270.610395222517, 280.154268134939, 295.113146283789, 
    294.462890625, 343.558789356902, 376.039397674819, 444.536544160588, 
    481.177986083193, 686.330412051292, 803.625015916513, 1105.41039175659, 
    1399.48492720246, 1566.7039057006, 1673.91447801922, 1748.97455969826, 
    1757.03263947287, 1755.01059494337, 1730.55762954994, 1736.08806986676, 
    1760.09711709766, 1772.7148009339, 1802.66884580957, 1794.94826907427, 
    1900.22801070059, 2028.62003798449, 2135.43335336864, 2316.9899777286, 
    2385.31292296583, 2409.11736498448, 2380.03235787507, 2284.42800706941, 
    2158.5470687266, 2191.85384798669, 2167.99719283008, 2063.80999937337, 
    1892.21538667506, 1756.30077066711, 2050.98300182278, 2510.84063534346, 
    3525.65638132679, 4065.89147763595, 4184.09344016234, 4192.9957203794, 
    4176.52040583629, 4204.15042602484, 4227.2770929791, 4230.91935744515, 
    4243.4189752448, 4240.94521383708, 4215.88550062088, 4115.15579899852, 
    4067.41075981297, 4005.65546266988, 3851.13561742809, 3747.3412891297, 
    3680.35342550049, 3614.87707237321, 3623.18115674463, 3657.55357676614, 
    3664.73094727074, 3703.27398523229, 3721.27612304688, 3701.27916458277, 
    3667.21740137341, 3635.79119209501, 3551.12385027012, 3490.81301528781, 
    3363.66758052085, 3243.5297077478, 3065.78548661781, 2837.61030619227, 
    2528.63566793852, 2175.85428202735, 1818.42089596691, 1387.81446009238, 
    1069.66775510836, 694.750688071408, 536.125258972534, 329.863553600147, 
    270.610395222517, 190, 190, 140, 160, 140, 150, 150, 160, 160, 170, 170, 
    170, 160, 150, 130, 110, 100, 90, 70, 60, 50, 50, 40, 40, 40, 40, 40, 40, 
    40, 40, 0, -0, -0, -0, -0, -0, -0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0 ;
}
