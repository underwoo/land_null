netcdf atmos_mosaicXland_mosaic {
dimensions:
	stringlen = 255 ;
	ncells = 5311 ;
	two = 2 ;
variables:
	char contact(stringlen) ;
		contact:standard_name = "grid_contact_spec" ;
		contact:contact_spec_version = "0.2" ;
		contact:contact_type = "exchange" ;
		contact:parent1_cell = "tile1_cell" ;
		contact:parent2_cell = "tile2_cell" ;
		contact:xgrid_area_field = "xgrid_area" ;
		contact:distant_to_parent1_centroid = "tile1_distance" ;
		contact:distant_to_parent2_centroid = "tile2_distance" ;
	int tile1_cell(ncells, two) ;
		tile1_cell:standard_name = "parent_cell_indices_in_mosaic1" ;
	int tile2_cell(ncells, two) ;
		tile2_cell:standard_name = "parent_cell_indices_in_mosaic2" ;
	double xgrid_area(ncells) ;
		xgrid_area:standard_name = "exchange_grid_area" ;
		xgrid_area:units = "m2" ;
	double tile1_distance(ncells, two) ;
		tile1_distance:standard_name = "distance_from_parent1_cell_centroid" ;
	double tile2_distance(ncells, two) ;
		tile2_distance:standard_name = "distance_from_parent2_cell_centroid" ;
data:

 contact = "atmos_mosaic:tile1::land_mosaic:tile1" ;

 tile1_cell =
  1, 1,
  2, 1,
  3, 1,
  4, 1,
  5, 1,
  6, 1,
  7, 1,
  8, 1,
  9, 1,
  10, 1,
  11, 1,
  12, 1,
  13, 1,
  14, 1,
  15, 1,
  16, 1,
  17, 1,
  18, 1,
  19, 1,
  20, 1,
  21, 1,
  22, 1,
  23, 1,
  24, 1,
  25, 1,
  26, 1,
  27, 1,
  28, 1,
  29, 1,
  30, 1,
  31, 1,
  32, 1,
  33, 1,
  34, 1,
  35, 1,
  36, 1,
  37, 1,
  38, 1,
  39, 1,
  40, 1,
  41, 1,
  42, 1,
  43, 1,
  44, 1,
  45, 1,
  46, 1,
  47, 1,
  48, 1,
  49, 1,
  50, 1,
  51, 1,
  52, 1,
  53, 1,
  54, 1,
  55, 1,
  56, 1,
  57, 1,
  58, 1,
  59, 1,
  60, 1,
  61, 1,
  62, 1,
  63, 1,
  64, 1,
  65, 1,
  66, 1,
  67, 1,
  68, 1,
  69, 1,
  70, 1,
  71, 1,
  72, 1,
  73, 1,
  74, 1,
  75, 1,
  76, 1,
  77, 1,
  78, 1,
  79, 1,
  80, 1,
  81, 1,
  82, 1,
  83, 1,
  84, 1,
  85, 1,
  86, 1,
  87, 1,
  88, 1,
  89, 1,
  90, 1,
  91, 1,
  92, 1,
  93, 1,
  94, 1,
  95, 1,
  96, 1,
  97, 1,
  98, 1,
  99, 1,
  100, 1,
  101, 1,
  102, 1,
  103, 1,
  104, 1,
  105, 1,
  106, 1,
  107, 1,
  108, 1,
  109, 1,
  110, 1,
  111, 1,
  112, 1,
  113, 1,
  114, 1,
  115, 1,
  116, 1,
  117, 1,
  118, 1,
  119, 1,
  120, 1,
  121, 1,
  122, 1,
  123, 1,
  124, 1,
  125, 1,
  126, 1,
  127, 1,
  128, 1,
  129, 1,
  130, 1,
  131, 1,
  132, 1,
  133, 1,
  134, 1,
  135, 1,
  136, 1,
  137, 1,
  138, 1,
  139, 1,
  140, 1,
  141, 1,
  142, 1,
  143, 1,
  144, 1,
  1, 2,
  2, 2,
  3, 2,
  4, 2,
  5, 2,
  6, 2,
  7, 2,
  8, 2,
  9, 2,
  10, 2,
  11, 2,
  12, 2,
  13, 2,
  14, 2,
  15, 2,
  16, 2,
  17, 2,
  18, 2,
  19, 2,
  20, 2,
  21, 2,
  22, 2,
  23, 2,
  24, 2,
  25, 2,
  26, 2,
  27, 2,
  28, 2,
  29, 2,
  30, 2,
  31, 2,
  32, 2,
  33, 2,
  34, 2,
  35, 2,
  36, 2,
  37, 2,
  38, 2,
  39, 2,
  40, 2,
  41, 2,
  42, 2,
  43, 2,
  44, 2,
  45, 2,
  46, 2,
  47, 2,
  48, 2,
  49, 2,
  50, 2,
  51, 2,
  52, 2,
  53, 2,
  54, 2,
  55, 2,
  56, 2,
  57, 2,
  58, 2,
  59, 2,
  60, 2,
  61, 2,
  62, 2,
  63, 2,
  64, 2,
  65, 2,
  66, 2,
  67, 2,
  68, 2,
  69, 2,
  70, 2,
  71, 2,
  72, 2,
  73, 2,
  74, 2,
  75, 2,
  76, 2,
  77, 2,
  78, 2,
  79, 2,
  80, 2,
  81, 2,
  82, 2,
  83, 2,
  84, 2,
  85, 2,
  86, 2,
  87, 2,
  88, 2,
  89, 2,
  90, 2,
  91, 2,
  92, 2,
  93, 2,
  94, 2,
  95, 2,
  96, 2,
  97, 2,
  98, 2,
  99, 2,
  100, 2,
  101, 2,
  102, 2,
  103, 2,
  104, 2,
  105, 2,
  106, 2,
  107, 2,
  108, 2,
  109, 2,
  110, 2,
  111, 2,
  112, 2,
  113, 2,
  114, 2,
  115, 2,
  116, 2,
  117, 2,
  118, 2,
  119, 2,
  120, 2,
  121, 2,
  122, 2,
  123, 2,
  124, 2,
  125, 2,
  126, 2,
  127, 2,
  128, 2,
  129, 2,
  130, 2,
  131, 2,
  132, 2,
  133, 2,
  134, 2,
  135, 2,
  136, 2,
  137, 2,
  138, 2,
  139, 2,
  140, 2,
  141, 2,
  142, 2,
  143, 2,
  144, 2,
  1, 3,
  2, 3,
  3, 3,
  4, 3,
  5, 3,
  6, 3,
  7, 3,
  8, 3,
  9, 3,
  10, 3,
  11, 3,
  12, 3,
  13, 3,
  14, 3,
  15, 3,
  16, 3,
  17, 3,
  18, 3,
  19, 3,
  20, 3,
  21, 3,
  22, 3,
  23, 3,
  24, 3,
  25, 3,
  26, 3,
  27, 3,
  28, 3,
  29, 3,
  30, 3,
  31, 3,
  32, 3,
  33, 3,
  34, 3,
  35, 3,
  36, 3,
  37, 3,
  38, 3,
  39, 3,
  40, 3,
  41, 3,
  42, 3,
  43, 3,
  44, 3,
  45, 3,
  46, 3,
  47, 3,
  48, 3,
  49, 3,
  50, 3,
  51, 3,
  52, 3,
  53, 3,
  54, 3,
  55, 3,
  56, 3,
  57, 3,
  58, 3,
  59, 3,
  60, 3,
  61, 3,
  62, 3,
  63, 3,
  64, 3,
  65, 3,
  66, 3,
  67, 3,
  68, 3,
  69, 3,
  70, 3,
  71, 3,
  72, 3,
  73, 3,
  74, 3,
  75, 3,
  76, 3,
  77, 3,
  78, 3,
  79, 3,
  80, 3,
  81, 3,
  82, 3,
  83, 3,
  84, 3,
  85, 3,
  86, 3,
  87, 3,
  88, 3,
  89, 3,
  90, 3,
  91, 3,
  92, 3,
  93, 3,
  94, 3,
  95, 3,
  96, 3,
  97, 3,
  98, 3,
  99, 3,
  100, 3,
  101, 3,
  102, 3,
  103, 3,
  104, 3,
  105, 3,
  106, 3,
  107, 3,
  108, 3,
  109, 3,
  110, 3,
  111, 3,
  112, 3,
  113, 3,
  114, 3,
  115, 3,
  116, 3,
  117, 3,
  118, 3,
  119, 3,
  120, 3,
  121, 3,
  122, 3,
  123, 3,
  124, 3,
  125, 3,
  126, 3,
  127, 3,
  128, 3,
  129, 3,
  130, 3,
  131, 3,
  132, 3,
  133, 3,
  134, 3,
  135, 3,
  136, 3,
  137, 3,
  138, 3,
  139, 3,
  140, 3,
  141, 3,
  142, 3,
  143, 3,
  144, 3,
  1, 4,
  2, 4,
  3, 4,
  4, 4,
  5, 4,
  6, 4,
  7, 4,
  8, 4,
  9, 4,
  10, 4,
  11, 4,
  12, 4,
  13, 4,
  14, 4,
  15, 4,
  16, 4,
  17, 4,
  18, 4,
  19, 4,
  20, 4,
  21, 4,
  22, 4,
  23, 4,
  24, 4,
  25, 4,
  26, 4,
  27, 4,
  28, 4,
  29, 4,
  30, 4,
  31, 4,
  32, 4,
  33, 4,
  34, 4,
  35, 4,
  36, 4,
  37, 4,
  38, 4,
  39, 4,
  40, 4,
  41, 4,
  42, 4,
  43, 4,
  44, 4,
  45, 4,
  46, 4,
  47, 4,
  48, 4,
  49, 4,
  50, 4,
  51, 4,
  52, 4,
  53, 4,
  54, 4,
  55, 4,
  56, 4,
  57, 4,
  58, 4,
  59, 4,
  60, 4,
  61, 4,
  62, 4,
  63, 4,
  64, 4,
  65, 4,
  66, 4,
  67, 4,
  68, 4,
  69, 4,
  70, 4,
  71, 4,
  72, 4,
  73, 4,
  74, 4,
  75, 4,
  76, 4,
  77, 4,
  78, 4,
  79, 4,
  80, 4,
  81, 4,
  82, 4,
  83, 4,
  84, 4,
  85, 4,
  86, 4,
  87, 4,
  88, 4,
  89, 4,
  90, 4,
  91, 4,
  92, 4,
  93, 4,
  94, 4,
  95, 4,
  96, 4,
  97, 4,
  98, 4,
  99, 4,
  100, 4,
  101, 4,
  102, 4,
  103, 4,
  104, 4,
  105, 4,
  106, 4,
  107, 4,
  108, 4,
  109, 4,
  110, 4,
  111, 4,
  112, 4,
  113, 4,
  114, 4,
  115, 4,
  116, 4,
  117, 4,
  118, 4,
  119, 4,
  120, 4,
  121, 4,
  122, 4,
  123, 4,
  124, 4,
  125, 4,
  126, 4,
  127, 4,
  128, 4,
  129, 4,
  130, 4,
  131, 4,
  132, 4,
  133, 4,
  134, 4,
  135, 4,
  136, 4,
  137, 4,
  138, 4,
  139, 4,
  140, 4,
  141, 4,
  142, 4,
  143, 4,
  144, 4,
  1, 5,
  2, 5,
  3, 5,
  4, 5,
  5, 5,
  6, 5,
  7, 5,
  8, 5,
  9, 5,
  10, 5,
  11, 5,
  12, 5,
  13, 5,
  14, 5,
  15, 5,
  16, 5,
  17, 5,
  18, 5,
  19, 5,
  20, 5,
  21, 5,
  22, 5,
  23, 5,
  24, 5,
  25, 5,
  26, 5,
  27, 5,
  28, 5,
  29, 5,
  30, 5,
  31, 5,
  32, 5,
  33, 5,
  34, 5,
  35, 5,
  36, 5,
  37, 5,
  38, 5,
  39, 5,
  40, 5,
  41, 5,
  42, 5,
  43, 5,
  44, 5,
  45, 5,
  46, 5,
  47, 5,
  48, 5,
  49, 5,
  50, 5,
  51, 5,
  52, 5,
  53, 5,
  54, 5,
  55, 5,
  56, 5,
  57, 5,
  58, 5,
  59, 5,
  60, 5,
  61, 5,
  62, 5,
  63, 5,
  64, 5,
  65, 5,
  66, 5,
  67, 5,
  68, 5,
  69, 5,
  70, 5,
  71, 5,
  72, 5,
  73, 5,
  74, 5,
  75, 5,
  76, 5,
  77, 5,
  78, 5,
  79, 5,
  80, 5,
  81, 5,
  82, 5,
  83, 5,
  84, 5,
  85, 5,
  86, 5,
  87, 5,
  88, 5,
  89, 5,
  90, 5,
  91, 5,
  92, 5,
  93, 5,
  94, 5,
  95, 5,
  96, 5,
  97, 5,
  98, 5,
  99, 5,
  100, 5,
  101, 5,
  102, 5,
  103, 5,
  104, 5,
  105, 5,
  106, 5,
  107, 5,
  108, 5,
  109, 5,
  110, 5,
  111, 5,
  112, 5,
  113, 5,
  114, 5,
  115, 5,
  116, 5,
  117, 5,
  118, 5,
  119, 5,
  120, 5,
  121, 5,
  122, 5,
  123, 5,
  124, 5,
  125, 5,
  126, 5,
  127, 5,
  128, 5,
  129, 5,
  130, 5,
  131, 5,
  132, 5,
  133, 5,
  134, 5,
  135, 5,
  136, 5,
  137, 5,
  138, 5,
  139, 5,
  140, 5,
  141, 5,
  142, 5,
  143, 5,
  144, 5,
  1, 6,
  2, 6,
  3, 6,
  4, 6,
  5, 6,
  6, 6,
  7, 6,
  8, 6,
  9, 6,
  10, 6,
  11, 6,
  12, 6,
  13, 6,
  14, 6,
  15, 6,
  16, 6,
  17, 6,
  18, 6,
  19, 6,
  20, 6,
  21, 6,
  22, 6,
  23, 6,
  24, 6,
  25, 6,
  26, 6,
  27, 6,
  28, 6,
  29, 6,
  30, 6,
  31, 6,
  32, 6,
  33, 6,
  34, 6,
  35, 6,
  36, 6,
  37, 6,
  38, 6,
  39, 6,
  40, 6,
  41, 6,
  42, 6,
  43, 6,
  44, 6,
  45, 6,
  46, 6,
  47, 6,
  48, 6,
  49, 6,
  50, 6,
  51, 6,
  52, 6,
  53, 6,
  54, 6,
  55, 6,
  56, 6,
  57, 6,
  58, 6,
  59, 6,
  60, 6,
  61, 6,
  62, 6,
  63, 6,
  64, 6,
  65, 6,
  66, 6,
  67, 6,
  68, 6,
  69, 6,
  70, 6,
  71, 6,
  72, 6,
  73, 6,
  74, 6,
  75, 6,
  76, 6,
  77, 6,
  78, 6,
  79, 6,
  80, 6,
  81, 6,
  82, 6,
  83, 6,
  84, 6,
  85, 6,
  86, 6,
  87, 6,
  88, 6,
  89, 6,
  90, 6,
  91, 6,
  92, 6,
  93, 6,
  94, 6,
  95, 6,
  96, 6,
  97, 6,
  98, 6,
  99, 6,
  100, 6,
  101, 6,
  102, 6,
  103, 6,
  104, 6,
  105, 6,
  106, 6,
  107, 6,
  108, 6,
  109, 6,
  110, 6,
  111, 6,
  112, 6,
  113, 6,
  114, 6,
  115, 6,
  116, 6,
  117, 6,
  118, 6,
  119, 6,
  120, 6,
  121, 6,
  122, 6,
  123, 6,
  124, 6,
  125, 6,
  126, 6,
  127, 6,
  128, 6,
  129, 6,
  130, 6,
  131, 6,
  132, 6,
  133, 6,
  134, 6,
  135, 6,
  136, 6,
  137, 6,
  138, 6,
  139, 6,
  140, 6,
  141, 6,
  142, 6,
  143, 6,
  144, 6,
  1, 7,
  2, 7,
  3, 7,
  4, 7,
  5, 7,
  6, 7,
  7, 7,
  8, 7,
  9, 7,
  10, 7,
  11, 7,
  12, 7,
  13, 7,
  14, 7,
  15, 7,
  16, 7,
  17, 7,
  18, 7,
  19, 7,
  20, 7,
  21, 7,
  22, 7,
  23, 7,
  24, 7,
  25, 7,
  26, 7,
  27, 7,
  28, 7,
  29, 7,
  30, 7,
  31, 7,
  32, 7,
  33, 7,
  34, 7,
  35, 7,
  36, 7,
  37, 7,
  38, 7,
  39, 7,
  40, 7,
  41, 7,
  42, 7,
  43, 7,
  44, 7,
  45, 7,
  46, 7,
  47, 7,
  48, 7,
  49, 7,
  50, 7,
  51, 7,
  52, 7,
  53, 7,
  54, 7,
  55, 7,
  56, 7,
  57, 7,
  58, 7,
  59, 7,
  60, 7,
  61, 7,
  62, 7,
  63, 7,
  64, 7,
  65, 7,
  66, 7,
  67, 7,
  68, 7,
  69, 7,
  70, 7,
  71, 7,
  72, 7,
  73, 7,
  74, 7,
  75, 7,
  76, 7,
  77, 7,
  78, 7,
  79, 7,
  80, 7,
  81, 7,
  82, 7,
  83, 7,
  84, 7,
  85, 7,
  86, 7,
  87, 7,
  88, 7,
  89, 7,
  90, 7,
  91, 7,
  92, 7,
  93, 7,
  94, 7,
  95, 7,
  96, 7,
  97, 7,
  98, 7,
  99, 7,
  100, 7,
  101, 7,
  102, 7,
  103, 7,
  104, 7,
  105, 7,
  106, 7,
  107, 7,
  108, 7,
  109, 7,
  110, 7,
  111, 7,
  112, 7,
  113, 7,
  114, 7,
  115, 7,
  116, 7,
  117, 7,
  118, 7,
  119, 7,
  120, 7,
  121, 7,
  122, 7,
  123, 7,
  124, 7,
  125, 7,
  126, 7,
  127, 7,
  128, 7,
  129, 7,
  130, 7,
  131, 7,
  132, 7,
  133, 7,
  134, 7,
  135, 7,
  136, 7,
  137, 7,
  138, 7,
  139, 7,
  140, 7,
  141, 7,
  142, 7,
  143, 7,
  144, 7,
  1, 8,
  2, 8,
  3, 8,
  4, 8,
  5, 8,
  6, 8,
  7, 8,
  8, 8,
  9, 8,
  10, 8,
  11, 8,
  12, 8,
  13, 8,
  14, 8,
  15, 8,
  16, 8,
  17, 8,
  18, 8,
  19, 8,
  20, 8,
  21, 8,
  22, 8,
  23, 8,
  24, 8,
  25, 8,
  26, 8,
  27, 8,
  28, 8,
  29, 8,
  30, 8,
  31, 8,
  32, 8,
  33, 8,
  34, 8,
  35, 8,
  36, 8,
  37, 8,
  38, 8,
  39, 8,
  40, 8,
  41, 8,
  42, 8,
  43, 8,
  44, 8,
  45, 8,
  46, 8,
  47, 8,
  48, 8,
  49, 8,
  50, 8,
  51, 8,
  52, 8,
  53, 8,
  54, 8,
  55, 8,
  56, 8,
  57, 8,
  58, 8,
  59, 8,
  60, 8,
  61, 8,
  62, 8,
  63, 8,
  64, 8,
  65, 8,
  66, 8,
  85, 8,
  86, 8,
  87, 8,
  88, 8,
  89, 8,
  90, 8,
  91, 8,
  92, 8,
  93, 8,
  94, 8,
  95, 8,
  96, 8,
  97, 8,
  98, 8,
  99, 8,
  100, 8,
  101, 8,
  102, 8,
  103, 8,
  104, 8,
  105, 8,
  106, 8,
  107, 8,
  108, 8,
  109, 8,
  110, 8,
  111, 8,
  112, 8,
  113, 8,
  114, 8,
  115, 8,
  116, 8,
  117, 8,
  118, 8,
  119, 8,
  120, 8,
  121, 8,
  122, 8,
  123, 8,
  133, 8,
  134, 8,
  135, 8,
  136, 8,
  137, 8,
  138, 8,
  139, 8,
  140, 8,
  141, 8,
  142, 8,
  143, 8,
  144, 8,
  1, 9,
  2, 9,
  3, 9,
  4, 9,
  5, 9,
  6, 9,
  7, 9,
  8, 9,
  9, 9,
  10, 9,
  11, 9,
  12, 9,
  13, 9,
  14, 9,
  15, 9,
  16, 9,
  17, 9,
  18, 9,
  19, 9,
  20, 9,
  21, 9,
  22, 9,
  23, 9,
  24, 9,
  25, 9,
  26, 9,
  27, 9,
  28, 9,
  29, 9,
  30, 9,
  31, 9,
  32, 9,
  33, 9,
  34, 9,
  35, 9,
  36, 9,
  37, 9,
  38, 9,
  39, 9,
  40, 9,
  41, 9,
  42, 9,
  43, 9,
  44, 9,
  45, 9,
  46, 9,
  47, 9,
  48, 9,
  49, 9,
  50, 9,
  51, 9,
  52, 9,
  53, 9,
  54, 9,
  55, 9,
  56, 9,
  57, 9,
  58, 9,
  59, 9,
  60, 9,
  61, 9,
  62, 9,
  63, 9,
  64, 9,
  65, 9,
  66, 9,
  67, 9,
  68, 9,
  91, 9,
  92, 9,
  93, 9,
  94, 9,
  95, 9,
  96, 9,
  97, 9,
  98, 9,
  99, 9,
  100, 9,
  101, 9,
  102, 9,
  103, 9,
  104, 9,
  105, 9,
  106, 9,
  107, 9,
  108, 9,
  109, 9,
  110, 9,
  111, 9,
  112, 9,
  113, 9,
  114, 9,
  115, 9,
  116, 9,
  117, 9,
  118, 9,
  119, 9,
  120, 9,
  121, 9,
  136, 9,
  137, 9,
  138, 9,
  139, 9,
  140, 9,
  141, 9,
  142, 9,
  143, 9,
  144, 9,
  1, 10,
  2, 10,
  3, 10,
  4, 10,
  5, 10,
  6, 10,
  7, 10,
  8, 10,
  9, 10,
  10, 10,
  11, 10,
  12, 10,
  13, 10,
  14, 10,
  15, 10,
  16, 10,
  17, 10,
  18, 10,
  19, 10,
  20, 10,
  21, 10,
  22, 10,
  23, 10,
  24, 10,
  25, 10,
  26, 10,
  27, 10,
  28, 10,
  29, 10,
  30, 10,
  31, 10,
  32, 10,
  33, 10,
  34, 10,
  35, 10,
  36, 10,
  37, 10,
  38, 10,
  39, 10,
  40, 10,
  41, 10,
  42, 10,
  43, 10,
  44, 10,
  45, 10,
  46, 10,
  47, 10,
  48, 10,
  49, 10,
  50, 10,
  51, 10,
  52, 10,
  53, 10,
  54, 10,
  55, 10,
  56, 10,
  57, 10,
  58, 10,
  59, 10,
  60, 10,
  61, 10,
  62, 10,
  63, 10,
  64, 10,
  65, 10,
  66, 10,
  67, 10,
  68, 10,
  69, 10,
  104, 10,
  105, 10,
  106, 10,
  107, 10,
  108, 10,
  113, 10,
  114, 10,
  115, 10,
  116, 10,
  117, 10,
  118, 10,
  119, 10,
  120, 10,
  138, 10,
  139, 10,
  140, 10,
  141, 10,
  142, 10,
  143, 10,
  144, 10,
  1, 11,
  2, 11,
  3, 11,
  4, 11,
  5, 11,
  6, 11,
  7, 11,
  8, 11,
  9, 11,
  10, 11,
  11, 11,
  12, 11,
  13, 11,
  14, 11,
  15, 11,
  16, 11,
  17, 11,
  18, 11,
  19, 11,
  20, 11,
  21, 11,
  22, 11,
  23, 11,
  24, 11,
  25, 11,
  26, 11,
  27, 11,
  28, 11,
  29, 11,
  30, 11,
  31, 11,
  32, 11,
  33, 11,
  34, 11,
  35, 11,
  36, 11,
  37, 11,
  38, 11,
  39, 11,
  40, 11,
  41, 11,
  42, 11,
  43, 11,
  44, 11,
  45, 11,
  46, 11,
  47, 11,
  48, 11,
  49, 11,
  50, 11,
  51, 11,
  52, 11,
  53, 11,
  54, 11,
  55, 11,
  56, 11,
  57, 11,
  58, 11,
  59, 11,
  60, 11,
  61, 11,
  62, 11,
  63, 11,
  64, 11,
  65, 11,
  66, 11,
  67, 11,
  114, 11,
  115, 11,
  116, 11,
  117, 11,
  118, 11,
  119, 11,
  120, 11,
  143, 11,
  144, 11,
  14, 12,
  17, 12,
  18, 12,
  19, 12,
  20, 12,
  21, 12,
  22, 12,
  23, 12,
  24, 12,
  25, 12,
  26, 12,
  27, 12,
  28, 12,
  32, 12,
  33, 12,
  34, 12,
  35, 12,
  36, 12,
  37, 12,
  38, 12,
  39, 12,
  40, 12,
  41, 12,
  42, 12,
  43, 12,
  44, 12,
  45, 12,
  46, 12,
  47, 12,
  48, 12,
  49, 12,
  50, 12,
  51, 12,
  52, 12,
  53, 12,
  54, 12,
  55, 12,
  56, 12,
  57, 12,
  58, 12,
  59, 12,
  60, 12,
  61, 12,
  62, 12,
  117, 12,
  118, 12,
  119, 12,
  120, 12,
  21, 13,
  22, 13,
  23, 13,
  35, 13,
  36, 13,
  38, 13,
  39, 13,
  40, 13,
  41, 13,
  42, 13,
  43, 13,
  44, 13,
  45, 13,
  46, 13,
  47, 13,
  51, 13,
  53, 13,
  54, 13,
  55, 13,
  56, 13,
  118, 13,
  119, 13,
  120, 13,
  121, 13,
  122, 13,
  119, 14,
  120, 14,
  121, 14,
  122, 14,
  115, 18,
  116, 18,
  117, 18,
  118, 18,
  115, 19,
  116, 19,
  117, 19,
  118, 19,
  114, 20,
  115, 20,
  116, 20,
  117, 20,
  120, 20,
  121, 20,
  28, 21,
  114, 21,
  115, 21,
  116, 21,
  117, 21,
  118, 21,
  68, 22,
  114, 22,
  115, 22,
  116, 22,
  117, 22,
  118, 22,
  67, 23,
  68, 23,
  69, 23,
  115, 23,
  116, 23,
  117, 23,
  118, 23,
  59, 24,
  60, 24,
  68, 24,
  69, 24,
  70, 24,
  115, 24,
  116, 24,
  117, 24,
  118, 24,
  59, 25,
  60, 25,
  69, 25,
  70, 25,
  71, 25,
  115, 25,
  116, 25,
  117, 25,
  118, 25,
  119, 25,
  120, 25,
  58, 26,
  59, 26,
  70, 26,
  71, 26,
  72, 26,
  115, 26,
  116, 26,
  117, 26,
  118, 26,
  119, 26,
  120, 26,
  121, 26,
  57, 27,
  58, 27,
  59, 27,
  60, 27,
  70, 27,
  71, 27,
  72, 27,
  115, 27,
  116, 27,
  117, 27,
  118, 27,
  119, 27,
  120, 27,
  121, 27,
  122, 27,
  47, 28,
  48, 28,
  55, 28,
  56, 28,
  57, 28,
  58, 28,
  59, 28,
  60, 28,
  61, 28,
  70, 28,
  115, 28,
  116, 28,
  117, 28,
  118, 28,
  119, 28,
  120, 28,
  121, 28,
  122, 28,
  123, 28,
  8, 29,
  9, 29,
  10, 29,
  11, 29,
  12, 29,
  47, 29,
  48, 29,
  49, 29,
  50, 29,
  51, 29,
  54, 29,
  55, 29,
  56, 29,
  57, 29,
  58, 29,
  59, 29,
  60, 29,
  61, 29,
  116, 29,
  117, 29,
  118, 29,
  119, 29,
  120, 29,
  121, 29,
  122, 29,
  123, 29,
  124, 29,
  7, 30,
  8, 30,
  9, 30,
  10, 30,
  11, 30,
  12, 30,
  13, 30,
  47, 30,
  48, 30,
  49, 30,
  50, 30,
  51, 30,
  52, 30,
  53, 30,
  54, 30,
  55, 30,
  56, 30,
  57, 30,
  58, 30,
  59, 30,
  60, 30,
  61, 30,
  62, 30,
  116, 30,
  117, 30,
  118, 30,
  119, 30,
  120, 30,
  121, 30,
  122, 30,
  123, 30,
  124, 30,
  7, 31,
  8, 31,
  9, 31,
  10, 31,
  11, 31,
  12, 31,
  13, 31,
  47, 31,
  48, 31,
  49, 31,
  50, 31,
  51, 31,
  52, 31,
  53, 31,
  54, 31,
  55, 31,
  56, 31,
  57, 31,
  58, 31,
  59, 31,
  60, 31,
  61, 31,
  62, 31,
  116, 31,
  117, 31,
  118, 31,
  119, 31,
  120, 31,
  121, 31,
  122, 31,
  123, 31,
  124, 31,
  125, 31,
  7, 32,
  8, 32,
  9, 32,
  10, 32,
  11, 32,
  12, 32,
  13, 32,
  14, 32,
  46, 32,
  47, 32,
  48, 32,
  49, 32,
  50, 32,
  51, 32,
  52, 32,
  53, 32,
  54, 32,
  55, 32,
  56, 32,
  57, 32,
  58, 32,
  59, 32,
  60, 32,
  61, 32,
  62, 32,
  116, 32,
  117, 32,
  118, 32,
  119, 32,
  120, 32,
  121, 32,
  122, 32,
  123, 32,
  124, 32,
  125, 32,
  7, 33,
  8, 33,
  9, 33,
  10, 33,
  11, 33,
  12, 33,
  13, 33,
  14, 33,
  18, 33,
  19, 33,
  46, 33,
  47, 33,
  48, 33,
  49, 33,
  50, 33,
  51, 33,
  52, 33,
  53, 33,
  54, 33,
  55, 33,
  56, 33,
  57, 33,
  58, 33,
  59, 33,
  60, 33,
  61, 33,
  62, 33,
  116, 33,
  117, 33,
  118, 33,
  119, 33,
  120, 33,
  121, 33,
  122, 33,
  123, 33,
  124, 33,
  125, 33,
  126, 33,
  6, 34,
  7, 34,
  8, 34,
  9, 34,
  10, 34,
  11, 34,
  12, 34,
  13, 34,
  14, 34,
  18, 34,
  19, 34,
  20, 34,
  46, 34,
  47, 34,
  48, 34,
  49, 34,
  50, 34,
  51, 34,
  52, 34,
  53, 34,
  54, 34,
  55, 34,
  56, 34,
  57, 34,
  58, 34,
  59, 34,
  60, 34,
  61, 34,
  116, 34,
  117, 34,
  118, 34,
  119, 34,
  120, 34,
  121, 34,
  122, 34,
  123, 34,
  124, 34,
  125, 34,
  126, 34,
  127, 34,
  128, 34,
  6, 35,
  7, 35,
  8, 35,
  9, 35,
  10, 35,
  11, 35,
  12, 35,
  13, 35,
  14, 35,
  18, 35,
  19, 35,
  20, 35,
  23, 35,
  46, 35,
  47, 35,
  48, 35,
  49, 35,
  50, 35,
  51, 35,
  52, 35,
  53, 35,
  54, 35,
  55, 35,
  56, 35,
  57, 35,
  58, 35,
  59, 35,
  60, 35,
  61, 35,
  67, 35,
  117, 35,
  118, 35,
  119, 35,
  120, 35,
  121, 35,
  122, 35,
  123, 35,
  124, 35,
  125, 35,
  126, 35,
  127, 35,
  128, 35,
  5, 36,
  6, 36,
  7, 36,
  8, 36,
  9, 36,
  10, 36,
  11, 36,
  12, 36,
  13, 36,
  14, 36,
  15, 36,
  18, 36,
  19, 36,
  20, 36,
  48, 36,
  49, 36,
  50, 36,
  51, 36,
  52, 36,
  53, 36,
  54, 36,
  55, 36,
  56, 36,
  57, 36,
  58, 36,
  59, 36,
  60, 36,
  117, 36,
  118, 36,
  119, 36,
  120, 36,
  121, 36,
  122, 36,
  123, 36,
  124, 36,
  125, 36,
  126, 36,
  127, 36,
  128, 36,
  5, 37,
  6, 37,
  7, 37,
  8, 37,
  9, 37,
  10, 37,
  11, 37,
  12, 37,
  13, 37,
  14, 37,
  15, 37,
  16, 37,
  18, 37,
  19, 37,
  20, 37,
  49, 37,
  50, 37,
  51, 37,
  52, 37,
  53, 37,
  54, 37,
  55, 37,
  56, 37,
  57, 37,
  58, 37,
  59, 37,
  71, 37,
  72, 37,
  115, 37,
  116, 37,
  117, 37,
  118, 37,
  119, 37,
  120, 37,
  121, 37,
  122, 37,
  123, 37,
  124, 37,
  125, 37,
  126, 37,
  127, 37,
  128, 37,
  129, 37,
  5, 38,
  6, 38,
  7, 38,
  8, 38,
  9, 38,
  10, 38,
  11, 38,
  12, 38,
  13, 38,
  14, 38,
  15, 38,
  16, 38,
  19, 38,
  20, 38,
  50, 38,
  51, 38,
  52, 38,
  53, 38,
  54, 38,
  55, 38,
  57, 38,
  58, 38,
  59, 38,
  114, 38,
  115, 38,
  116, 38,
  117, 38,
  118, 38,
  119, 38,
  120, 38,
  121, 38,
  122, 38,
  123, 38,
  124, 38,
  125, 38,
  126, 38,
  127, 38,
  128, 38,
  129, 38,
  5, 39,
  6, 39,
  7, 39,
  8, 39,
  9, 39,
  10, 39,
  11, 39,
  12, 39,
  13, 39,
  14, 39,
  15, 39,
  16, 39,
  20, 39,
  51, 39,
  52, 39,
  53, 39,
  54, 39,
  55, 39,
  57, 39,
  58, 39,
  114, 39,
  115, 39,
  116, 39,
  117, 39,
  118, 39,
  119, 39,
  120, 39,
  121, 39,
  122, 39,
  123, 39,
  124, 39,
  125, 39,
  126, 39,
  127, 39,
  128, 39,
  129, 39,
  6, 40,
  7, 40,
  8, 40,
  9, 40,
  10, 40,
  11, 40,
  12, 40,
  13, 40,
  14, 40,
  15, 40,
  16, 40,
  50, 40,
  53, 40,
  54, 40,
  55, 40,
  57, 40,
  58, 40,
  61, 40,
  113, 40,
  114, 40,
  115, 40,
  116, 40,
  117, 40,
  118, 40,
  119, 40,
  120, 40,
  121, 40,
  122, 40,
  123, 40,
  124, 40,
  125, 40,
  126, 40,
  127, 40,
  128, 40,
  129, 40,
  130, 40,
  6, 41,
  7, 41,
  8, 41,
  9, 41,
  10, 41,
  11, 41,
  12, 41,
  13, 41,
  14, 41,
  15, 41,
  16, 41,
  47, 41,
  48, 41,
  49, 41,
  50, 41,
  51, 41,
  57, 41,
  58, 41,
  59, 41,
  60, 41,
  61, 41,
  113, 41,
  114, 41,
  115, 41,
  116, 41,
  117, 41,
  118, 41,
  119, 41,
  120, 41,
  121, 41,
  122, 41,
  123, 41,
  124, 41,
  125, 41,
  126, 41,
  127, 41,
  128, 41,
  129, 41,
  130, 41,
  5, 42,
  6, 42,
  7, 42,
  8, 42,
  9, 42,
  10, 42,
  11, 42,
  12, 42,
  13, 42,
  14, 42,
  15, 42,
  16, 42,
  43, 42,
  44, 42,
  45, 42,
  46, 42,
  47, 42,
  48, 42,
  49, 42,
  53, 42,
  54, 42,
  56, 42,
  57, 42,
  58, 42,
  59, 42,
  60, 42,
  61, 42,
  63, 42,
  112, 42,
  113, 42,
  114, 42,
  115, 42,
  116, 42,
  117, 42,
  118, 42,
  119, 42,
  120, 42,
  121, 42,
  122, 42,
  123, 42,
  124, 42,
  125, 42,
  126, 42,
  127, 42,
  128, 42,
  129, 42,
  130, 42,
  5, 43,
  6, 43,
  7, 43,
  8, 43,
  9, 43,
  10, 43,
  11, 43,
  12, 43,
  13, 43,
  14, 43,
  15, 43,
  16, 43,
  41, 43,
  42, 43,
  43, 43,
  48, 43,
  49, 43,
  50, 43,
  54, 43,
  55, 43,
  56, 43,
  57, 43,
  58, 43,
  59, 43,
  60, 43,
  61, 43,
  112, 43,
  113, 43,
  114, 43,
  115, 43,
  116, 43,
  117, 43,
  118, 43,
  119, 43,
  120, 43,
  121, 43,
  122, 43,
  123, 43,
  124, 43,
  125, 43,
  126, 43,
  127, 43,
  128, 43,
  129, 43,
  130, 43,
  4, 44,
  5, 44,
  6, 44,
  7, 44,
  8, 44,
  9, 44,
  10, 44,
  11, 44,
  12, 44,
  13, 44,
  14, 44,
  15, 44,
  16, 44,
  17, 44,
  41, 44,
  42, 44,
  43, 44,
  45, 44,
  46, 44,
  47, 44,
  48, 44,
  49, 44,
  50, 44,
  51, 44,
  52, 44,
  53, 44,
  54, 44,
  55, 44,
  56, 44,
  57, 44,
  58, 44,
  112, 44,
  113, 44,
  114, 44,
  115, 44,
  116, 44,
  117, 44,
  118, 44,
  119, 44,
  120, 44,
  121, 44,
  122, 44,
  123, 44,
  124, 44,
  125, 44,
  126, 44,
  127, 44,
  128, 44,
  129, 44,
  4, 45,
  5, 45,
  6, 45,
  7, 45,
  8, 45,
  9, 45,
  10, 45,
  11, 45,
  12, 45,
  13, 45,
  14, 45,
  15, 45,
  16, 45,
  17, 45,
  18, 45,
  41, 45,
  42, 45,
  43, 45,
  44, 45,
  45, 45,
  46, 45,
  47, 45,
  48, 45,
  49, 45,
  50, 45,
  51, 45,
  52, 45,
  53, 45,
  54, 45,
  55, 45,
  56, 45,
  112, 45,
  113, 45,
  114, 45,
  115, 45,
  116, 45,
  117, 45,
  118, 45,
  119, 45,
  120, 45,
  121, 45,
  122, 45,
  123, 45,
  124, 45,
  125, 45,
  126, 45,
  4, 46,
  5, 46,
  6, 46,
  7, 46,
  8, 46,
  9, 46,
  10, 46,
  11, 46,
  12, 46,
  13, 46,
  14, 46,
  15, 46,
  16, 46,
  17, 46,
  18, 46,
  39, 46,
  40, 46,
  41, 46,
  42, 46,
  44, 46,
  45, 46,
  46, 46,
  47, 46,
  48, 46,
  49, 46,
  50, 46,
  51, 46,
  52, 46,
  113, 46,
  114, 46,
  115, 46,
  116, 46,
  117, 46,
  118, 46,
  119, 46,
  120, 46,
  121, 46,
  122, 46,
  123, 46,
  124, 46,
  4, 47,
  5, 47,
  6, 47,
  7, 47,
  8, 47,
  9, 47,
  10, 47,
  11, 47,
  12, 47,
  13, 47,
  14, 47,
  15, 47,
  16, 47,
  17, 47,
  18, 47,
  19, 47,
  20, 47,
  39, 47,
  40, 47,
  41, 47,
  42, 47,
  44, 47,
  45, 47,
  46, 47,
  47, 47,
  48, 47,
  52, 47,
  113, 47,
  114, 47,
  115, 47,
  116, 47,
  117, 47,
  118, 47,
  119, 47,
  120, 47,
  121, 47,
  122, 47,
  123, 47,
  124, 47,
  1, 48,
  3, 48,
  4, 48,
  5, 48,
  6, 48,
  7, 48,
  8, 48,
  9, 48,
  10, 48,
  11, 48,
  12, 48,
  13, 48,
  14, 48,
  15, 48,
  16, 48,
  17, 48,
  18, 48,
  19, 48,
  20, 48,
  39, 48,
  40, 48,
  41, 48,
  42, 48,
  46, 48,
  47, 48,
  48, 48,
  51, 48,
  114, 48,
  115, 48,
  116, 48,
  117, 48,
  118, 48,
  119, 48,
  120, 48,
  121, 48,
  122, 48,
  123, 48,
  124, 48,
  141, 48,
  142, 48,
  143, 48,
  144, 48,
  1, 49,
  2, 49,
  3, 49,
  4, 49,
  5, 49,
  6, 49,
  7, 49,
  8, 49,
  9, 49,
  10, 49,
  11, 49,
  12, 49,
  13, 49,
  14, 49,
  15, 49,
  16, 49,
  17, 49,
  18, 49,
  19, 49,
  20, 49,
  31, 49,
  32, 49,
  33, 49,
  40, 49,
  41, 49,
  42, 49,
  47, 49,
  48, 49,
  49, 49,
  50, 49,
  51, 49,
  111, 49,
  112, 49,
  113, 49,
  114, 49,
  115, 49,
  116, 49,
  117, 49,
  118, 49,
  119, 49,
  120, 49,
  121, 49,
  122, 49,
  139, 49,
  140, 49,
  141, 49,
  142, 49,
  143, 49,
  144, 49,
  1, 50,
  2, 50,
  3, 50,
  4, 50,
  5, 50,
  6, 50,
  7, 50,
  8, 50,
  9, 50,
  10, 50,
  11, 50,
  12, 50,
  13, 50,
  14, 50,
  15, 50,
  16, 50,
  17, 50,
  18, 50,
  19, 50,
  20, 50,
  21, 50,
  31, 50,
  32, 50,
  33, 50,
  40, 50,
  42, 50,
  43, 50,
  44, 50,
  47, 50,
  48, 50,
  50, 50,
  51, 50,
  110, 50,
  111, 50,
  112, 50,
  113, 50,
  114, 50,
  115, 50,
  116, 50,
  117, 50,
  118, 50,
  119, 50,
  120, 50,
  139, 50,
  140, 50,
  141, 50,
  142, 50,
  143, 50,
  144, 50,
  1, 51,
  2, 51,
  3, 51,
  4, 51,
  5, 51,
  6, 51,
  7, 51,
  8, 51,
  9, 51,
  10, 51,
  11, 51,
  12, 51,
  13, 51,
  14, 51,
  15, 51,
  16, 51,
  17, 51,
  18, 51,
  19, 51,
  20, 51,
  21, 51,
  31, 51,
  32, 51,
  40, 51,
  41, 51,
  42, 51,
  43, 51,
  44, 51,
  48, 51,
  49, 51,
  50, 51,
  110, 51,
  111, 51,
  115, 51,
  116, 51,
  117, 51,
  118, 51,
  119, 51,
  120, 51,
  138, 51,
  139, 51,
  140, 51,
  141, 51,
  142, 51,
  143, 51,
  144, 51,
  1, 52,
  2, 52,
  3, 52,
  4, 52,
  5, 52,
  6, 52,
  7, 52,
  8, 52,
  9, 52,
  10, 52,
  11, 52,
  12, 52,
  13, 52,
  14, 52,
  15, 52,
  16, 52,
  17, 52,
  18, 52,
  19, 52,
  20, 52,
  30, 52,
  31, 52,
  32, 52,
  40, 52,
  41, 52,
  42, 52,
  43, 52,
  44, 52,
  49, 52,
  50, 52,
  108, 52,
  109, 52,
  110, 52,
  111, 52,
  138, 52,
  139, 52,
  140, 52,
  141, 52,
  142, 52,
  143, 52,
  144, 52,
  1, 53,
  2, 53,
  3, 53,
  4, 53,
  5, 53,
  6, 53,
  7, 53,
  8, 53,
  9, 53,
  10, 53,
  11, 53,
  12, 53,
  13, 53,
  14, 53,
  15, 53,
  16, 53,
  17, 53,
  18, 53,
  19, 53,
  20, 53,
  21, 53,
  30, 53,
  31, 53,
  32, 53,
  33, 53,
  40, 53,
  41, 53,
  42, 53,
  43, 53,
  44, 53,
  49, 53,
  105, 53,
  106, 53,
  107, 53,
  108, 53,
  109, 53,
  110, 53,
  111, 53,
  138, 53,
  139, 53,
  140, 53,
  141, 53,
  142, 53,
  143, 53,
  144, 53,
  1, 54,
  2, 54,
  3, 54,
  4, 54,
  5, 54,
  6, 54,
  7, 54,
  8, 54,
  9, 54,
  10, 54,
  11, 54,
  12, 54,
  13, 54,
  14, 54,
  15, 54,
  16, 54,
  17, 54,
  18, 54,
  19, 54,
  20, 54,
  21, 54,
  22, 54,
  23, 54,
  30, 54,
  31, 54,
  32, 54,
  33, 54,
  34, 54,
  38, 54,
  39, 54,
  40, 54,
  41, 54,
  42, 54,
  43, 54,
  44, 54,
  49, 54,
  103, 54,
  104, 54,
  105, 54,
  106, 54,
  107, 54,
  108, 54,
  109, 54,
  115, 54,
  116, 54,
  118, 54,
  138, 54,
  139, 54,
  140, 54,
  141, 54,
  142, 54,
  143, 54,
  144, 54,
  1, 55,
  2, 55,
  3, 55,
  4, 55,
  5, 55,
  6, 55,
  7, 55,
  8, 55,
  9, 55,
  10, 55,
  11, 55,
  12, 55,
  13, 55,
  14, 55,
  15, 55,
  16, 55,
  17, 55,
  18, 55,
  19, 55,
  20, 55,
  21, 55,
  22, 55,
  23, 55,
  24, 55,
  30, 55,
  31, 55,
  32, 55,
  33, 55,
  34, 55,
  35, 55,
  38, 55,
  39, 55,
  40, 55,
  41, 55,
  42, 55,
  43, 55,
  44, 55,
  45, 55,
  82, 55,
  103, 55,
  104, 55,
  105, 55,
  106, 55,
  108, 55,
  109, 55,
  114, 55,
  115, 55,
  116, 55,
  117, 55,
  118, 55,
  138, 55,
  139, 55,
  140, 55,
  141, 55,
  142, 55,
  143, 55,
  144, 55,
  1, 56,
  2, 56,
  3, 56,
  4, 56,
  5, 56,
  6, 56,
  7, 56,
  8, 56,
  9, 56,
  10, 56,
  11, 56,
  12, 56,
  13, 56,
  14, 56,
  15, 56,
  16, 56,
  17, 56,
  18, 56,
  19, 56,
  20, 56,
  21, 56,
  22, 56,
  23, 56,
  24, 56,
  28, 56,
  29, 56,
  30, 56,
  31, 56,
  32, 56,
  33, 56,
  34, 56,
  35, 56,
  36, 56,
  37, 56,
  38, 56,
  39, 56,
  40, 56,
  41, 56,
  42, 56,
  43, 56,
  44, 56,
  45, 56,
  46, 56,
  49, 56,
  82, 56,
  102, 56,
  103, 56,
  104, 56,
  105, 56,
  106, 56,
  109, 56,
  111, 56,
  112, 56,
  113, 56,
  114, 56,
  138, 56,
  139, 56,
  140, 56,
  141, 56,
  142, 56,
  143, 56,
  144, 56,
  1, 57,
  2, 57,
  3, 57,
  4, 57,
  5, 57,
  6, 57,
  7, 57,
  8, 57,
  9, 57,
  10, 57,
  11, 57,
  12, 57,
  13, 57,
  14, 57,
  15, 57,
  16, 57,
  17, 57,
  18, 57,
  19, 57,
  20, 57,
  21, 57,
  22, 57,
  23, 57,
  24, 57,
  27, 57,
  28, 57,
  29, 57,
  30, 57,
  31, 57,
  32, 57,
  33, 57,
  34, 57,
  35, 57,
  36, 57,
  37, 57,
  38, 57,
  39, 57,
  40, 57,
  41, 57,
  42, 57,
  43, 57,
  44, 57,
  45, 57,
  46, 57,
  47, 57,
  48, 57,
  49, 57,
  100, 57,
  101, 57,
  102, 57,
  103, 57,
  104, 57,
  105, 57,
  111, 57,
  112, 57,
  113, 57,
  138, 57,
  139, 57,
  140, 57,
  141, 57,
  142, 57,
  143, 57,
  144, 57,
  1, 58,
  2, 58,
  3, 58,
  4, 58,
  5, 58,
  6, 58,
  7, 58,
  8, 58,
  9, 58,
  10, 58,
  11, 58,
  12, 58,
  13, 58,
  14, 58,
  15, 58,
  16, 58,
  17, 58,
  18, 58,
  19, 58,
  20, 58,
  21, 58,
  22, 58,
  23, 58,
  24, 58,
  25, 58,
  26, 58,
  27, 58,
  28, 58,
  29, 58,
  30, 58,
  31, 58,
  32, 58,
  33, 58,
  34, 58,
  35, 58,
  36, 58,
  37, 58,
  38, 58,
  39, 58,
  40, 58,
  41, 58,
  42, 58,
  43, 58,
  44, 58,
  45, 58,
  46, 58,
  47, 58,
  48, 58,
  49, 58,
  99, 58,
  100, 58,
  101, 58,
  102, 58,
  103, 58,
  104, 58,
  105, 58,
  106, 58,
  112, 58,
  139, 58,
  140, 58,
  141, 58,
  142, 58,
  143, 58,
  144, 58,
  1, 59,
  2, 59,
  3, 59,
  4, 59,
  5, 59,
  6, 59,
  7, 59,
  8, 59,
  9, 59,
  10, 59,
  11, 59,
  12, 59,
  13, 59,
  14, 59,
  15, 59,
  16, 59,
  17, 59,
  18, 59,
  19, 59,
  20, 59,
  21, 59,
  22, 59,
  23, 59,
  24, 59,
  25, 59,
  26, 59,
  27, 59,
  28, 59,
  29, 59,
  30, 59,
  31, 59,
  32, 59,
  33, 59,
  34, 59,
  35, 59,
  36, 59,
  37, 59,
  38, 59,
  39, 59,
  40, 59,
  41, 59,
  42, 59,
  43, 59,
  44, 59,
  45, 59,
  46, 59,
  47, 59,
  48, 59,
  49, 59,
  99, 59,
  100, 59,
  101, 59,
  102, 59,
  103, 59,
  104, 59,
  105, 59,
  106, 59,
  111, 59,
  112, 59,
  139, 59,
  140, 59,
  141, 59,
  142, 59,
  143, 59,
  144, 59,
  1, 60,
  2, 60,
  3, 60,
  4, 60,
  5, 60,
  6, 60,
  7, 60,
  8, 60,
  9, 60,
  10, 60,
  11, 60,
  12, 60,
  13, 60,
  14, 60,
  15, 60,
  16, 60,
  17, 60,
  18, 60,
  19, 60,
  20, 60,
  21, 60,
  22, 60,
  23, 60,
  24, 60,
  25, 60,
  26, 60,
  27, 60,
  28, 60,
  29, 60,
  30, 60,
  31, 60,
  32, 60,
  33, 60,
  34, 60,
  35, 60,
  36, 60,
  37, 60,
  38, 60,
  39, 60,
  40, 60,
  41, 60,
  42, 60,
  43, 60,
  44, 60,
  45, 60,
  46, 60,
  47, 60,
  48, 60,
  49, 60,
  98, 60,
  99, 60,
  100, 60,
  101, 60,
  102, 60,
  103, 60,
  104, 60,
  105, 60,
  106, 60,
  107, 60,
  108, 60,
  109, 60,
  110, 60,
  111, 60,
  112, 60,
  140, 60,
  141, 60,
  142, 60,
  143, 60,
  144, 60,
  1, 61,
  2, 61,
  3, 61,
  4, 61,
  5, 61,
  6, 61,
  7, 61,
  8, 61,
  9, 61,
  10, 61,
  11, 61,
  12, 61,
  13, 61,
  14, 61,
  15, 61,
  16, 61,
  17, 61,
  18, 61,
  19, 61,
  20, 61,
  21, 61,
  22, 61,
  23, 61,
  24, 61,
  25, 61,
  26, 61,
  27, 61,
  28, 61,
  29, 61,
  30, 61,
  31, 61,
  32, 61,
  33, 61,
  34, 61,
  35, 61,
  36, 61,
  37, 61,
  38, 61,
  39, 61,
  40, 61,
  41, 61,
  42, 61,
  43, 61,
  44, 61,
  45, 61,
  46, 61,
  47, 61,
  48, 61,
  49, 61,
  53, 61,
  98, 61,
  99, 61,
  100, 61,
  101, 61,
  102, 61,
  103, 61,
  104, 61,
  105, 61,
  106, 61,
  107, 61,
  108, 61,
  109, 61,
  110, 61,
  111, 61,
  112, 61,
  141, 61,
  142, 61,
  143, 61,
  144, 61,
  1, 62,
  2, 62,
  3, 62,
  4, 62,
  5, 62,
  6, 62,
  9, 62,
  10, 62,
  15, 62,
  16, 62,
  17, 62,
  18, 62,
  19, 62,
  20, 62,
  21, 62,
  22, 62,
  23, 62,
  24, 62,
  25, 62,
  26, 62,
  27, 62,
  28, 62,
  29, 62,
  30, 62,
  31, 62,
  32, 62,
  33, 62,
  34, 62,
  35, 62,
  36, 62,
  37, 62,
  38, 62,
  39, 62,
  40, 62,
  41, 62,
  42, 62,
  43, 62,
  44, 62,
  45, 62,
  46, 62,
  47, 62,
  48, 62,
  49, 62,
  51, 62,
  53, 62,
  54, 62,
  55, 62,
  97, 62,
  98, 62,
  99, 62,
  100, 62,
  101, 62,
  102, 62,
  103, 62,
  104, 62,
  105, 62,
  106, 62,
  107, 62,
  108, 62,
  109, 62,
  110, 62,
  111, 62,
  112, 62,
  113, 62,
  114, 62,
  141, 62,
  142, 62,
  143, 62,
  144, 62,
  1, 63,
  2, 63,
  3, 63,
  4, 63,
  5, 63,
  12, 63,
  13, 63,
  14, 63,
  15, 63,
  16, 63,
  17, 63,
  18, 63,
  19, 63,
  20, 63,
  21, 63,
  22, 63,
  23, 63,
  24, 63,
  25, 63,
  26, 63,
  27, 63,
  28, 63,
  29, 63,
  30, 63,
  31, 63,
  32, 63,
  33, 63,
  34, 63,
  35, 63,
  36, 63,
  37, 63,
  38, 63,
  39, 63,
  40, 63,
  41, 63,
  42, 63,
  43, 63,
  44, 63,
  45, 63,
  46, 63,
  47, 63,
  48, 63,
  49, 63,
  51, 63,
  52, 63,
  53, 63,
  54, 63,
  55, 63,
  56, 63,
  57, 63,
  96, 63,
  97, 63,
  98, 63,
  99, 63,
  100, 63,
  101, 63,
  102, 63,
  103, 63,
  104, 63,
  105, 63,
  106, 63,
  107, 63,
  108, 63,
  109, 63,
  110, 63,
  111, 63,
  112, 63,
  113, 63,
  114, 63,
  142, 63,
  143, 63,
  144, 63,
  1, 64,
  2, 64,
  3, 64,
  4, 64,
  5, 64,
  6, 64,
  7, 64,
  9, 64,
  10, 64,
  11, 64,
  12, 64,
  13, 64,
  14, 64,
  15, 64,
  16, 64,
  17, 64,
  18, 64,
  19, 64,
  20, 64,
  21, 64,
  22, 64,
  23, 64,
  24, 64,
  25, 64,
  26, 64,
  27, 64,
  28, 64,
  29, 64,
  30, 64,
  31, 64,
  32, 64,
  33, 64,
  34, 64,
  35, 64,
  36, 64,
  37, 64,
  38, 64,
  39, 64,
  40, 64,
  41, 64,
  42, 64,
  43, 64,
  44, 64,
  45, 64,
  46, 64,
  47, 64,
  48, 64,
  49, 64,
  51, 64,
  52, 64,
  55, 64,
  56, 64,
  57, 64,
  95, 64,
  96, 64,
  97, 64,
  98, 64,
  99, 64,
  100, 64,
  101, 64,
  102, 64,
  103, 64,
  104, 64,
  105, 64,
  106, 64,
  107, 64,
  108, 64,
  109, 64,
  110, 64,
  111, 64,
  112, 64,
  113, 64,
  114, 64,
  141, 64,
  142, 64,
  143, 64,
  144, 64,
  1, 65,
  4, 65,
  6, 65,
  7, 65,
  8, 65,
  9, 65,
  10, 65,
  11, 65,
  12, 65,
  13, 65,
  14, 65,
  15, 65,
  16, 65,
  17, 65,
  18, 65,
  19, 65,
  20, 65,
  21, 65,
  22, 65,
  23, 65,
  24, 65,
  25, 65,
  26, 65,
  27, 65,
  28, 65,
  29, 65,
  30, 65,
  31, 65,
  32, 65,
  33, 65,
  34, 65,
  35, 65,
  36, 65,
  37, 65,
  38, 65,
  39, 65,
  40, 65,
  41, 65,
  42, 65,
  43, 65,
  44, 65,
  45, 65,
  46, 65,
  47, 65,
  48, 65,
  49, 65,
  50, 65,
  51, 65,
  52, 65,
  56, 65,
  57, 65,
  95, 65,
  96, 65,
  97, 65,
  98, 65,
  99, 65,
  100, 65,
  101, 65,
  102, 65,
  103, 65,
  104, 65,
  105, 65,
  106, 65,
  107, 65,
  108, 65,
  109, 65,
  110, 65,
  111, 65,
  112, 65,
  113, 65,
  114, 65,
  115, 65,
  141, 65,
  142, 65,
  143, 65,
  144, 65,
  1, 66,
  2, 66,
  4, 66,
  5, 66,
  6, 66,
  7, 66,
  8, 66,
  9, 66,
  10, 66,
  11, 66,
  12, 66,
  13, 66,
  14, 66,
  15, 66,
  16, 66,
  17, 66,
  18, 66,
  19, 66,
  20, 66,
  21, 66,
  22, 66,
  23, 66,
  24, 66,
  25, 66,
  26, 66,
  27, 66,
  28, 66,
  29, 66,
  30, 66,
  31, 66,
  32, 66,
  33, 66,
  34, 66,
  35, 66,
  36, 66,
  37, 66,
  38, 66,
  39, 66,
  40, 66,
  41, 66,
  42, 66,
  43, 66,
  44, 66,
  45, 66,
  46, 66,
  47, 66,
  48, 66,
  49, 66,
  50, 66,
  51, 66,
  52, 66,
  53, 66,
  57, 66,
  58, 66,
  95, 66,
  96, 66,
  97, 66,
  98, 66,
  99, 66,
  100, 66,
  101, 66,
  102, 66,
  103, 66,
  104, 66,
  105, 66,
  106, 66,
  107, 66,
  108, 66,
  109, 66,
  110, 66,
  111, 66,
  112, 66,
  113, 66,
  114, 66,
  115, 66,
  116, 66,
  141, 66,
  142, 66,
  143, 66,
  144, 66,
  1, 67,
  2, 67,
  3, 67,
  4, 67,
  5, 67,
  6, 67,
  7, 67,
  8, 67,
  9, 67,
  10, 67,
  11, 67,
  12, 67,
  16, 67,
  17, 67,
  18, 67,
  19, 67,
  20, 67,
  21, 67,
  22, 67,
  23, 67,
  24, 67,
  25, 67,
  26, 67,
  27, 67,
  28, 67,
  29, 67,
  30, 67,
  31, 67,
  32, 67,
  33, 67,
  34, 67,
  35, 67,
  36, 67,
  37, 67,
  38, 67,
  39, 67,
  40, 67,
  41, 67,
  42, 67,
  43, 67,
  44, 67,
  45, 67,
  46, 67,
  47, 67,
  48, 67,
  49, 67,
  50, 67,
  51, 67,
  52, 67,
  53, 67,
  54, 67,
  55, 67,
  57, 67,
  58, 67,
  95, 67,
  96, 67,
  97, 67,
  98, 67,
  99, 67,
  100, 67,
  101, 67,
  102, 67,
  103, 67,
  104, 67,
  105, 67,
  106, 67,
  107, 67,
  108, 67,
  109, 67,
  110, 67,
  111, 67,
  112, 67,
  113, 67,
  114, 67,
  115, 67,
  116, 67,
  117, 67,
  118, 67,
  119, 67,
  141, 67,
  142, 67,
  143, 67,
  144, 67,
  1, 68,
  2, 68,
  3, 68,
  4, 68,
  5, 68,
  6, 68,
  7, 68,
  8, 68,
  9, 68,
  10, 68,
  11, 68,
  12, 68,
  13, 68,
  14, 68,
  15, 68,
  16, 68,
  17, 68,
  18, 68,
  19, 68,
  20, 68,
  21, 68,
  22, 68,
  23, 68,
  24, 68,
  25, 68,
  26, 68,
  27, 68,
  28, 68,
  29, 68,
  30, 68,
  31, 68,
  32, 68,
  33, 68,
  34, 68,
  35, 68,
  36, 68,
  37, 68,
  38, 68,
  39, 68,
  40, 68,
  41, 68,
  42, 68,
  43, 68,
  44, 68,
  45, 68,
  46, 68,
  47, 68,
  48, 68,
  49, 68,
  50, 68,
  51, 68,
  52, 68,
  53, 68,
  54, 68,
  55, 68,
  56, 68,
  57, 68,
  58, 68,
  95, 68,
  96, 68,
  97, 68,
  98, 68,
  99, 68,
  100, 68,
  101, 68,
  102, 68,
  103, 68,
  104, 68,
  105, 68,
  106, 68,
  107, 68,
  108, 68,
  109, 68,
  110, 68,
  111, 68,
  112, 68,
  113, 68,
  114, 68,
  115, 68,
  116, 68,
  117, 68,
  118, 68,
  119, 68,
  120, 68,
  144, 68,
  1, 69,
  2, 69,
  3, 69,
  4, 69,
  5, 69,
  6, 69,
  7, 69,
  8, 69,
  9, 69,
  10, 69,
  11, 69,
  12, 69,
  13, 69,
  14, 69,
  15, 69,
  16, 69,
  17, 69,
  18, 69,
  19, 69,
  20, 69,
  21, 69,
  22, 69,
  23, 69,
  24, 69,
  25, 69,
  26, 69,
  27, 69,
  28, 69,
  29, 69,
  30, 69,
  31, 69,
  32, 69,
  33, 69,
  34, 69,
  35, 69,
  36, 69,
  37, 69,
  38, 69,
  39, 69,
  40, 69,
  41, 69,
  42, 69,
  43, 69,
  44, 69,
  45, 69,
  46, 69,
  47, 69,
  48, 69,
  49, 69,
  50, 69,
  51, 69,
  52, 69,
  53, 69,
  54, 69,
  55, 69,
  56, 69,
  57, 69,
  58, 69,
  95, 69,
  96, 69,
  97, 69,
  98, 69,
  99, 69,
  100, 69,
  101, 69,
  102, 69,
  103, 69,
  104, 69,
  105, 69,
  106, 69,
  107, 69,
  108, 69,
  109, 69,
  110, 69,
  111, 69,
  112, 69,
  113, 69,
  114, 69,
  115, 69,
  116, 69,
  117, 69,
  118, 69,
  119, 69,
  121, 69,
  122, 69,
  123, 69,
  143, 69,
  144, 69,
  1, 70,
  2, 70,
  3, 70,
  4, 70,
  5, 70,
  6, 70,
  7, 70,
  8, 70,
  9, 70,
  10, 70,
  11, 70,
  12, 70,
  13, 70,
  14, 70,
  15, 70,
  16, 70,
  17, 70,
  18, 70,
  19, 70,
  20, 70,
  21, 70,
  22, 70,
  23, 70,
  24, 70,
  25, 70,
  26, 70,
  27, 70,
  28, 70,
  29, 70,
  30, 70,
  31, 70,
  32, 70,
  33, 70,
  34, 70,
  35, 70,
  36, 70,
  37, 70,
  38, 70,
  39, 70,
  40, 70,
  41, 70,
  42, 70,
  43, 70,
  44, 70,
  45, 70,
  46, 70,
  47, 70,
  48, 70,
  49, 70,
  50, 70,
  51, 70,
  52, 70,
  53, 70,
  54, 70,
  55, 70,
  56, 70,
  57, 70,
  58, 70,
  93, 70,
  94, 70,
  95, 70,
  96, 70,
  97, 70,
  98, 70,
  99, 70,
  100, 70,
  101, 70,
  102, 70,
  103, 70,
  104, 70,
  105, 70,
  106, 70,
  107, 70,
  108, 70,
  109, 70,
  110, 70,
  111, 70,
  112, 70,
  113, 70,
  114, 70,
  115, 70,
  116, 70,
  117, 70,
  118, 70,
  119, 70,
  120, 70,
  121, 70,
  122, 70,
  123, 70,
  143, 70,
  144, 70,
  1, 71,
  2, 71,
  3, 71,
  4, 71,
  5, 71,
  6, 71,
  7, 71,
  8, 71,
  9, 71,
  10, 71,
  11, 71,
  12, 71,
  13, 71,
  14, 71,
  15, 71,
  16, 71,
  17, 71,
  18, 71,
  19, 71,
  20, 71,
  21, 71,
  22, 71,
  23, 71,
  24, 71,
  25, 71,
  26, 71,
  27, 71,
  28, 71,
  29, 71,
  30, 71,
  31, 71,
  32, 71,
  33, 71,
  34, 71,
  35, 71,
  36, 71,
  37, 71,
  38, 71,
  39, 71,
  40, 71,
  41, 71,
  42, 71,
  43, 71,
  44, 71,
  45, 71,
  46, 71,
  47, 71,
  48, 71,
  49, 71,
  50, 71,
  51, 71,
  52, 71,
  53, 71,
  54, 71,
  55, 71,
  56, 71,
  57, 71,
  58, 71,
  63, 71,
  64, 71,
  93, 71,
  94, 71,
  95, 71,
  96, 71,
  97, 71,
  98, 71,
  99, 71,
  100, 71,
  101, 71,
  102, 71,
  103, 71,
  104, 71,
  105, 71,
  106, 71,
  107, 71,
  108, 71,
  109, 71,
  110, 71,
  111, 71,
  112, 71,
  113, 71,
  114, 71,
  115, 71,
  116, 71,
  117, 71,
  118, 71,
  119, 71,
  120, 71,
  121, 71,
  122, 71,
  141, 71,
  142, 71,
  143, 71,
  144, 71,
  1, 72,
  3, 72,
  4, 72,
  5, 72,
  6, 72,
  7, 72,
  8, 72,
  9, 72,
  10, 72,
  11, 72,
  12, 72,
  13, 72,
  14, 72,
  15, 72,
  16, 72,
  17, 72,
  18, 72,
  19, 72,
  20, 72,
  21, 72,
  22, 72,
  23, 72,
  24, 72,
  25, 72,
  26, 72,
  27, 72,
  28, 72,
  29, 72,
  30, 72,
  31, 72,
  32, 72,
  33, 72,
  34, 72,
  35, 72,
  36, 72,
  37, 72,
  38, 72,
  39, 72,
  40, 72,
  41, 72,
  42, 72,
  43, 72,
  44, 72,
  45, 72,
  46, 72,
  47, 72,
  48, 72,
  49, 72,
  50, 72,
  51, 72,
  52, 72,
  53, 72,
  54, 72,
  55, 72,
  56, 72,
  57, 72,
  58, 72,
  63, 72,
  64, 72,
  65, 72,
  77, 72,
  79, 72,
  92, 72,
  93, 72,
  94, 72,
  95, 72,
  96, 72,
  97, 72,
  98, 72,
  99, 72,
  100, 72,
  101, 72,
  102, 72,
  103, 72,
  104, 72,
  105, 72,
  106, 72,
  107, 72,
  108, 72,
  109, 72,
  110, 72,
  111, 72,
  112, 72,
  113, 72,
  114, 72,
  115, 72,
  116, 72,
  117, 72,
  118, 72,
  119, 72,
  120, 72,
  121, 72,
  122, 72,
  141, 72,
  142, 72,
  143, 72,
  144, 72,
  4, 73,
  5, 73,
  6, 73,
  7, 73,
  8, 73,
  9, 73,
  10, 73,
  11, 73,
  12, 73,
  13, 73,
  14, 73,
  15, 73,
  16, 73,
  17, 73,
  18, 73,
  19, 73,
  20, 73,
  21, 73,
  22, 73,
  23, 73,
  24, 73,
  25, 73,
  26, 73,
  27, 73,
  28, 73,
  29, 73,
  30, 73,
  31, 73,
  32, 73,
  33, 73,
  34, 73,
  35, 73,
  36, 73,
  37, 73,
  38, 73,
  39, 73,
  40, 73,
  41, 73,
  42, 73,
  43, 73,
  44, 73,
  45, 73,
  46, 73,
  47, 73,
  48, 73,
  49, 73,
  50, 73,
  51, 73,
  52, 73,
  53, 73,
  54, 73,
  55, 73,
  56, 73,
  63, 73,
  64, 73,
  65, 73,
  66, 73,
  79, 73,
  80, 73,
  81, 73,
  91, 73,
  92, 73,
  93, 73,
  94, 73,
  95, 73,
  96, 73,
  97, 73,
  98, 73,
  99, 73,
  100, 73,
  101, 73,
  102, 73,
  103, 73,
  104, 73,
  105, 73,
  106, 73,
  107, 73,
  108, 73,
  109, 73,
  110, 73,
  111, 73,
  112, 73,
  113, 73,
  114, 73,
  115, 73,
  116, 73,
  117, 73,
  118, 73,
  119, 73,
  120, 73,
  121, 73,
  122, 73,
  141, 73,
  142, 73,
  143, 73,
  144, 73,
  3, 74,
  4, 74,
  5, 74,
  6, 74,
  7, 74,
  9, 74,
  10, 74,
  11, 74,
  12, 74,
  13, 74,
  14, 74,
  15, 74,
  16, 74,
  17, 74,
  18, 74,
  19, 74,
  20, 74,
  21, 74,
  22, 74,
  23, 74,
  24, 74,
  25, 74,
  26, 74,
  27, 74,
  28, 74,
  29, 74,
  30, 74,
  31, 74,
  32, 74,
  33, 74,
  34, 74,
  35, 74,
  36, 74,
  37, 74,
  38, 74,
  39, 74,
  40, 74,
  41, 74,
  42, 74,
  43, 74,
  44, 74,
  45, 74,
  46, 74,
  47, 74,
  48, 74,
  49, 74,
  50, 74,
  51, 74,
  52, 74,
  53, 74,
  54, 74,
  55, 74,
  56, 74,
  57, 74,
  63, 74,
  64, 74,
  65, 74,
  66, 74,
  80, 74,
  81, 74,
  82, 74,
  83, 74,
  84, 74,
  89, 74,
  90, 74,
  91, 74,
  92, 74,
  93, 74,
  94, 74,
  95, 74,
  96, 74,
  97, 74,
  98, 74,
  99, 74,
  100, 74,
  101, 74,
  102, 74,
  103, 74,
  104, 74,
  105, 74,
  106, 74,
  107, 74,
  108, 74,
  109, 74,
  113, 74,
  114, 74,
  115, 74,
  116, 74,
  117, 74,
  118, 74,
  119, 74,
  120, 74,
  142, 74,
  143, 74,
  144, 74,
  3, 75,
  4, 75,
  5, 75,
  6, 75,
  7, 75,
  8, 75,
  9, 75,
  10, 75,
  11, 75,
  12, 75,
  13, 75,
  14, 75,
  15, 75,
  16, 75,
  17, 75,
  18, 75,
  19, 75,
  20, 75,
  21, 75,
  22, 75,
  23, 75,
  24, 75,
  25, 75,
  26, 75,
  27, 75,
  28, 75,
  29, 75,
  30, 75,
  31, 75,
  32, 75,
  33, 75,
  34, 75,
  35, 75,
  36, 75,
  37, 75,
  38, 75,
  39, 75,
  40, 75,
  41, 75,
  42, 75,
  43, 75,
  44, 75,
  45, 75,
  46, 75,
  47, 75,
  48, 75,
  49, 75,
  50, 75,
  51, 75,
  52, 75,
  53, 75,
  54, 75,
  55, 75,
  56, 75,
  57, 75,
  58, 75,
  59, 75,
  60, 75,
  61, 75,
  62, 75,
  64, 75,
  65, 75,
  66, 75,
  67, 75,
  68, 75,
  69, 75,
  78, 75,
  79, 75,
  80, 75,
  81, 75,
  82, 75,
  83, 75,
  84, 75,
  85, 75,
  86, 75,
  87, 75,
  88, 75,
  89, 75,
  90, 75,
  91, 75,
  92, 75,
  93, 75,
  94, 75,
  95, 75,
  96, 75,
  97, 75,
  98, 75,
  99, 75,
  100, 75,
  101, 75,
  102, 75,
  103, 75,
  104, 75,
  105, 75,
  106, 75,
  107, 75,
  113, 75,
  114, 75,
  115, 75,
  116, 75,
  117, 75,
  118, 75,
  119, 75,
  126, 75,
  127, 75,
  143, 75,
  144, 75,
  3, 76,
  4, 76,
  5, 76,
  6, 76,
  7, 76,
  8, 76,
  9, 76,
  10, 76,
  11, 76,
  12, 76,
  13, 76,
  14, 76,
  15, 76,
  16, 76,
  17, 76,
  18, 76,
  19, 76,
  20, 76,
  21, 76,
  22, 76,
  23, 76,
  24, 76,
  25, 76,
  26, 76,
  27, 76,
  28, 76,
  29, 76,
  30, 76,
  31, 76,
  32, 76,
  33, 76,
  34, 76,
  35, 76,
  36, 76,
  37, 76,
  38, 76,
  39, 76,
  40, 76,
  41, 76,
  42, 76,
  43, 76,
  44, 76,
  45, 76,
  46, 76,
  47, 76,
  48, 76,
  49, 76,
  50, 76,
  51, 76,
  52, 76,
  53, 76,
  54, 76,
  55, 76,
  56, 76,
  57, 76,
  58, 76,
  59, 76,
  60, 76,
  61, 76,
  62, 76,
  63, 76,
  64, 76,
  65, 76,
  66, 76,
  67, 76,
  68, 76,
  69, 76,
  70, 76,
  71, 76,
  72, 76,
  78, 76,
  79, 76,
  80, 76,
  81, 76,
  82, 76,
  83, 76,
  84, 76,
  85, 76,
  86, 76,
  87, 76,
  88, 76,
  89, 76,
  90, 76,
  91, 76,
  92, 76,
  93, 76,
  94, 76,
  95, 76,
  96, 76,
  97, 76,
  98, 76,
  99, 76,
  100, 76,
  101, 76,
  102, 76,
  103, 76,
  104, 76,
  105, 76,
  106, 76,
  107, 76,
  108, 76,
  113, 76,
  114, 76,
  115, 76,
  116, 76,
  117, 76,
  118, 76,
  125, 76,
  126, 76,
  127, 76,
  128, 76,
  141, 76,
  142, 76,
  144, 76,
  3, 77,
  4, 77,
  5, 77,
  6, 77,
  7, 77,
  8, 77,
  9, 77,
  10, 77,
  11, 77,
  12, 77,
  13, 77,
  14, 77,
  15, 77,
  16, 77,
  17, 77,
  18, 77,
  19, 77,
  20, 77,
  21, 77,
  22, 77,
  23, 77,
  24, 77,
  25, 77,
  26, 77,
  27, 77,
  28, 77,
  29, 77,
  30, 77,
  31, 77,
  32, 77,
  33, 77,
  34, 77,
  35, 77,
  36, 77,
  37, 77,
  38, 77,
  39, 77,
  40, 77,
  41, 77,
  42, 77,
  43, 77,
  44, 77,
  45, 77,
  46, 77,
  47, 77,
  48, 77,
  49, 77,
  50, 77,
  51, 77,
  52, 77,
  53, 77,
  54, 77,
  55, 77,
  56, 77,
  57, 77,
  58, 77,
  59, 77,
  60, 77,
  61, 77,
  62, 77,
  63, 77,
  64, 77,
  65, 77,
  66, 77,
  67, 77,
  68, 77,
  69, 77,
  70, 77,
  71, 77,
  72, 77,
  75, 77,
  76, 77,
  78, 77,
  79, 77,
  80, 77,
  81, 77,
  82, 77,
  83, 77,
  84, 77,
  85, 77,
  86, 77,
  87, 77,
  88, 77,
  89, 77,
  90, 77,
  91, 77,
  92, 77,
  93, 77,
  94, 77,
  95, 77,
  96, 77,
  97, 77,
  98, 77,
  99, 77,
  100, 77,
  101, 77,
  102, 77,
  103, 77,
  104, 77,
  105, 77,
  106, 77,
  107, 77,
  108, 77,
  109, 77,
  110, 77,
  111, 77,
  112, 77,
  113, 77,
  114, 77,
  115, 77,
  116, 77,
  117, 77,
  118, 77,
  119, 77,
  124, 77,
  125, 77,
  126, 77,
  127, 77,
  128, 77,
  136, 77,
  137, 77,
  138, 77,
  139, 77,
  141, 77,
  142, 77,
  5, 78,
  6, 78,
  7, 78,
  8, 78,
  9, 78,
  10, 78,
  11, 78,
  12, 78,
  13, 78,
  14, 78,
  15, 78,
  16, 78,
  17, 78,
  18, 78,
  19, 78,
  20, 78,
  21, 78,
  22, 78,
  23, 78,
  24, 78,
  25, 78,
  26, 78,
  27, 78,
  28, 78,
  29, 78,
  30, 78,
  31, 78,
  32, 78,
  33, 78,
  34, 78,
  35, 78,
  36, 78,
  37, 78,
  38, 78,
  39, 78,
  40, 78,
  41, 78,
  42, 78,
  43, 78,
  44, 78,
  45, 78,
  46, 78,
  47, 78,
  48, 78,
  49, 78,
  50, 78,
  51, 78,
  52, 78,
  53, 78,
  54, 78,
  55, 78,
  56, 78,
  57, 78,
  58, 78,
  59, 78,
  60, 78,
  61, 78,
  62, 78,
  63, 78,
  64, 78,
  65, 78,
  66, 78,
  67, 78,
  68, 78,
  69, 78,
  70, 78,
  71, 78,
  72, 78,
  73, 78,
  74, 78,
  75, 78,
  76, 78,
  77, 78,
  78, 78,
  79, 78,
  80, 78,
  81, 78,
  82, 78,
  83, 78,
  84, 78,
  85, 78,
  86, 78,
  87, 78,
  88, 78,
  89, 78,
  90, 78,
  91, 78,
  92, 78,
  93, 78,
  94, 78,
  95, 78,
  96, 78,
  97, 78,
  98, 78,
  99, 78,
  100, 78,
  101, 78,
  102, 78,
  103, 78,
  104, 78,
  105, 78,
  106, 78,
  107, 78,
  108, 78,
  109, 78,
  110, 78,
  111, 78,
  112, 78,
  113, 78,
  114, 78,
  115, 78,
  116, 78,
  117, 78,
  118, 78,
  119, 78,
  120, 78,
  123, 78,
  124, 78,
  125, 78,
  126, 78,
  127, 78,
  128, 78,
  129, 78,
  130, 78,
  131, 78,
  135, 78,
  136, 78,
  137, 78,
  138, 78,
  139, 78,
  6, 79,
  7, 79,
  8, 79,
  9, 79,
  10, 79,
  11, 79,
  12, 79,
  13, 79,
  14, 79,
  15, 79,
  16, 79,
  17, 79,
  18, 79,
  19, 79,
  20, 79,
  21, 79,
  22, 79,
  23, 79,
  24, 79,
  25, 79,
  26, 79,
  27, 79,
  28, 79,
  29, 79,
  30, 79,
  31, 79,
  32, 79,
  33, 79,
  34, 79,
  35, 79,
  36, 79,
  37, 79,
  38, 79,
  39, 79,
  40, 79,
  41, 79,
  42, 79,
  43, 79,
  44, 79,
  45, 79,
  46, 79,
  47, 79,
  48, 79,
  49, 79,
  50, 79,
  51, 79,
  52, 79,
  53, 79,
  54, 79,
  55, 79,
  56, 79,
  57, 79,
  58, 79,
  59, 79,
  60, 79,
  61, 79,
  62, 79,
  63, 79,
  64, 79,
  65, 79,
  66, 79,
  67, 79,
  68, 79,
  69, 79,
  70, 79,
  71, 79,
  72, 79,
  73, 79,
  74, 79,
  75, 79,
  76, 79,
  78, 79,
  79, 79,
  80, 79,
  81, 79,
  82, 79,
  83, 79,
  84, 79,
  85, 79,
  86, 79,
  87, 79,
  88, 79,
  89, 79,
  90, 79,
  91, 79,
  92, 79,
  93, 79,
  94, 79,
  95, 79,
  96, 79,
  97, 79,
  98, 79,
  99, 79,
  100, 79,
  101, 79,
  102, 79,
  103, 79,
  104, 79,
  105, 79,
  106, 79,
  107, 79,
  108, 79,
  109, 79,
  110, 79,
  111, 79,
  112, 79,
  114, 79,
  115, 79,
  116, 79,
  117, 79,
  118, 79,
  119, 79,
  120, 79,
  123, 79,
  124, 79,
  125, 79,
  126, 79,
  127, 79,
  128, 79,
  129, 79,
  130, 79,
  131, 79,
  132, 79,
  7, 80,
  8, 80,
  9, 80,
  10, 80,
  11, 80,
  12, 80,
  13, 80,
  14, 80,
  15, 80,
  16, 80,
  19, 80,
  20, 80,
  21, 80,
  22, 80,
  23, 80,
  24, 80,
  25, 80,
  26, 80,
  27, 80,
  28, 80,
  29, 80,
  30, 80,
  31, 80,
  32, 80,
  33, 80,
  34, 80,
  35, 80,
  36, 80,
  37, 80,
  38, 80,
  39, 80,
  40, 80,
  41, 80,
  42, 80,
  43, 80,
  44, 80,
  45, 80,
  46, 80,
  47, 80,
  48, 80,
  49, 80,
  50, 80,
  51, 80,
  52, 80,
  53, 80,
  54, 80,
  55, 80,
  56, 80,
  57, 80,
  58, 80,
  59, 80,
  60, 80,
  61, 80,
  62, 80,
  63, 80,
  64, 80,
  65, 80,
  66, 80,
  67, 80,
  68, 80,
  69, 80,
  70, 80,
  71, 80,
  72, 80,
  73, 80,
  78, 80,
  79, 80,
  80, 80,
  81, 80,
  82, 80,
  83, 80,
  84, 80,
  85, 80,
  86, 80,
  87, 80,
  88, 80,
  89, 80,
  90, 80,
  91, 80,
  92, 80,
  93, 80,
  94, 80,
  95, 80,
  96, 80,
  97, 80,
  98, 80,
  99, 80,
  100, 80,
  101, 80,
  102, 80,
  103, 80,
  104, 80,
  105, 80,
  106, 80,
  107, 80,
  108, 80,
  109, 80,
  110, 80,
  111, 80,
  112, 80,
  113, 80,
  114, 80,
  115, 80,
  116, 80,
  117, 80,
  118, 80,
  123, 80,
  124, 80,
  125, 80,
  126, 80,
  127, 80,
  128, 80,
  129, 80,
  130, 80,
  131, 80,
  132, 80,
  133, 80,
  134, 80,
  135, 80,
  9, 81,
  10, 81,
  11, 81,
  21, 81,
  22, 81,
  23, 81,
  27, 81,
  28, 81,
  29, 81,
  30, 81,
  31, 81,
  32, 81,
  33, 81,
  34, 81,
  35, 81,
  36, 81,
  37, 81,
  38, 81,
  39, 81,
  40, 81,
  41, 81,
  42, 81,
  43, 81,
  44, 81,
  45, 81,
  46, 81,
  47, 81,
  48, 81,
  49, 81,
  50, 81,
  51, 81,
  52, 81,
  53, 81,
  54, 81,
  55, 81,
  56, 81,
  57, 81,
  58, 81,
  59, 81,
  60, 81,
  61, 81,
  62, 81,
  63, 81,
  64, 81,
  72, 81,
  73, 81,
  81, 81,
  82, 81,
  83, 81,
  94, 81,
  95, 81,
  96, 81,
  97, 81,
  98, 81,
  99, 81,
  100, 81,
  101, 81,
  102, 81,
  103, 81,
  104, 81,
  105, 81,
  106, 81,
  107, 81,
  108, 81,
  109, 81,
  110, 81,
  111, 81,
  112, 81,
  113, 81,
  114, 81,
  115, 81,
  116, 81,
  117, 81,
  122, 81,
  123, 81,
  124, 81,
  125, 81,
  126, 81,
  127, 81,
  128, 81,
  129, 81,
  130, 81,
  131, 81,
  132, 81,
  133, 81,
  134, 81,
  135, 81,
  136, 81,
  21, 82,
  22, 82,
  23, 82,
  24, 82,
  28, 82,
  29, 82,
  30, 82,
  31, 82,
  32, 82,
  33, 82,
  34, 82,
  35, 82,
  36, 82,
  37, 82,
  38, 82,
  39, 82,
  40, 82,
  41, 82,
  42, 82,
  43, 82,
  44, 82,
  45, 82,
  46, 82,
  47, 82,
  48, 82,
  49, 82,
  50, 82,
  51, 82,
  52, 82,
  56, 82,
  57, 82,
  58, 82,
  59, 82,
  60, 82,
  61, 82,
  94, 82,
  95, 82,
  96, 82,
  97, 82,
  98, 82,
  99, 82,
  100, 82,
  101, 82,
  102, 82,
  103, 82,
  104, 82,
  105, 82,
  106, 82,
  107, 82,
  108, 82,
  109, 82,
  110, 82,
  111, 82,
  112, 82,
  113, 82,
  114, 82,
  122, 82,
  123, 82,
  124, 82,
  125, 82,
  126, 82,
  127, 82,
  128, 82,
  129, 82,
  130, 82,
  131, 82,
  132, 82,
  133, 82,
  134, 82,
  135, 82,
  136, 82,
  22, 83,
  23, 83,
  24, 83,
  25, 83,
  26, 83,
  27, 83,
  28, 83,
  35, 83,
  36, 83,
  37, 83,
  38, 83,
  39, 83,
  40, 83,
  41, 83,
  42, 83,
  43, 83,
  44, 83,
  45, 83,
  46, 83,
  47, 83,
  55, 83,
  56, 83,
  57, 83,
  58, 83,
  59, 83,
  60, 83,
  61, 83,
  95, 83,
  96, 83,
  97, 83,
  98, 83,
  99, 83,
  100, 83,
  101, 83,
  102, 83,
  103, 83,
  104, 83,
  105, 83,
  106, 83,
  107, 83,
  108, 83,
  109, 83,
  110, 83,
  111, 83,
  112, 83,
  113, 83,
  117, 83,
  118, 83,
  119, 83,
  120, 83,
  121, 83,
  122, 83,
  123, 83,
  124, 83,
  125, 83,
  126, 83,
  127, 83,
  128, 83,
  129, 83,
  130, 83,
  131, 83,
  132, 83,
  133, 83,
  134, 83,
  135, 83,
  136, 83,
  137, 83,
  5, 84,
  6, 84,
  7, 84,
  8, 84,
  9, 84,
  10, 84,
  26, 84,
  27, 84,
  39, 84,
  40, 84,
  41, 84,
  42, 84,
  43, 84,
  44, 84,
  45, 84,
  96, 84,
  97, 84,
  98, 84,
  99, 84,
  103, 84,
  104, 84,
  105, 84,
  106, 84,
  107, 84,
  108, 84,
  109, 84,
  110, 84,
  111, 84,
  112, 84,
  113, 84,
  114, 84,
  116, 84,
  117, 84,
  118, 84,
  119, 84,
  120, 84,
  121, 84,
  122, 84,
  123, 84,
  124, 84,
  125, 84,
  126, 84,
  127, 84,
  128, 84,
  129, 84,
  130, 84,
  131, 84,
  132, 84,
  133, 84,
  134, 84,
  135, 84,
  136, 84,
  137, 84,
  5, 85,
  6, 85,
  7, 85,
  8, 85,
  9, 85,
  10, 85,
  11, 85,
  12, 85,
  19, 85,
  20, 85,
  21, 85,
  22, 85,
  23, 85,
  24, 85,
  25, 85,
  26, 85,
  36, 85,
  37, 85,
  38, 85,
  39, 85,
  40, 85,
  41, 85,
  42, 85,
  43, 85,
  103, 85,
  104, 85,
  105, 85,
  106, 85,
  107, 85,
  108, 85,
  109, 85,
  110, 85,
  111, 85,
  112, 85,
  113, 85,
  114, 85,
  115, 85,
  116, 85,
  118, 85,
  119, 85,
  120, 85,
  121, 85,
  122, 85,
  123, 85,
  124, 85,
  125, 85,
  126, 85,
  127, 85,
  128, 85,
  129, 85,
  130, 85,
  131, 85,
  132, 85,
  133, 85,
  134, 85,
  135, 85,
  136, 85,
  137, 85,
  138, 85,
  20, 86,
  21, 86,
  22, 86,
  23, 86,
  25, 86,
  26, 86,
  37, 86,
  38, 86,
  39, 86,
  40, 86,
  107, 86,
  108, 86,
  109, 86,
  110, 86,
  111, 86,
  112, 86,
  113, 86,
  114, 86,
  115, 86,
  116, 86,
  117, 86,
  119, 86,
  120, 86,
  121, 86,
  122, 86,
  123, 86,
  124, 86,
  125, 86,
  126, 86,
  127, 86,
  128, 86,
  129, 86,
  130, 86,
  131, 86,
  132, 86,
  133, 86,
  134, 86,
  135, 86,
  136, 86,
  137, 86,
  138, 86,
  139, 86,
  111, 87,
  112, 87,
  113, 87,
  114, 87,
  115, 87,
  116, 87,
  117, 87,
  118, 87,
  127, 87,
  128, 87,
  129, 87,
  130, 87,
  131, 87,
  132, 87,
  133, 87,
  134, 87 ;

 tile2_cell =
  1, 1,
  2, 1,
  3, 1,
  4, 1,
  5, 1,
  6, 1,
  7, 1,
  8, 1,
  9, 1,
  10, 1,
  11, 1,
  12, 1,
  13, 1,
  14, 1,
  15, 1,
  16, 1,
  17, 1,
  18, 1,
  19, 1,
  20, 1,
  21, 1,
  22, 1,
  23, 1,
  24, 1,
  25, 1,
  26, 1,
  27, 1,
  28, 1,
  29, 1,
  30, 1,
  31, 1,
  32, 1,
  33, 1,
  34, 1,
  35, 1,
  36, 1,
  37, 1,
  38, 1,
  39, 1,
  40, 1,
  41, 1,
  42, 1,
  43, 1,
  44, 1,
  45, 1,
  46, 1,
  47, 1,
  48, 1,
  49, 1,
  50, 1,
  51, 1,
  52, 1,
  53, 1,
  54, 1,
  55, 1,
  56, 1,
  57, 1,
  58, 1,
  59, 1,
  60, 1,
  61, 1,
  62, 1,
  63, 1,
  64, 1,
  65, 1,
  66, 1,
  67, 1,
  68, 1,
  69, 1,
  70, 1,
  71, 1,
  72, 1,
  73, 1,
  74, 1,
  75, 1,
  76, 1,
  77, 1,
  78, 1,
  79, 1,
  80, 1,
  81, 1,
  82, 1,
  83, 1,
  84, 1,
  85, 1,
  86, 1,
  87, 1,
  88, 1,
  89, 1,
  90, 1,
  91, 1,
  92, 1,
  93, 1,
  94, 1,
  95, 1,
  96, 1,
  97, 1,
  98, 1,
  99, 1,
  100, 1,
  101, 1,
  102, 1,
  103, 1,
  104, 1,
  105, 1,
  106, 1,
  107, 1,
  108, 1,
  109, 1,
  110, 1,
  111, 1,
  112, 1,
  113, 1,
  114, 1,
  115, 1,
  116, 1,
  117, 1,
  118, 1,
  119, 1,
  120, 1,
  121, 1,
  122, 1,
  123, 1,
  124, 1,
  125, 1,
  126, 1,
  127, 1,
  128, 1,
  129, 1,
  130, 1,
  131, 1,
  132, 1,
  133, 1,
  134, 1,
  135, 1,
  136, 1,
  137, 1,
  138, 1,
  139, 1,
  140, 1,
  141, 1,
  142, 1,
  143, 1,
  144, 1,
  1, 2,
  2, 2,
  3, 2,
  4, 2,
  5, 2,
  6, 2,
  7, 2,
  8, 2,
  9, 2,
  10, 2,
  11, 2,
  12, 2,
  13, 2,
  14, 2,
  15, 2,
  16, 2,
  17, 2,
  18, 2,
  19, 2,
  20, 2,
  21, 2,
  22, 2,
  23, 2,
  24, 2,
  25, 2,
  26, 2,
  27, 2,
  28, 2,
  29, 2,
  30, 2,
  31, 2,
  32, 2,
  33, 2,
  34, 2,
  35, 2,
  36, 2,
  37, 2,
  38, 2,
  39, 2,
  40, 2,
  41, 2,
  42, 2,
  43, 2,
  44, 2,
  45, 2,
  46, 2,
  47, 2,
  48, 2,
  49, 2,
  50, 2,
  51, 2,
  52, 2,
  53, 2,
  54, 2,
  55, 2,
  56, 2,
  57, 2,
  58, 2,
  59, 2,
  60, 2,
  61, 2,
  62, 2,
  63, 2,
  64, 2,
  65, 2,
  66, 2,
  67, 2,
  68, 2,
  69, 2,
  70, 2,
  71, 2,
  72, 2,
  73, 2,
  74, 2,
  75, 2,
  76, 2,
  77, 2,
  78, 2,
  79, 2,
  80, 2,
  81, 2,
  82, 2,
  83, 2,
  84, 2,
  85, 2,
  86, 2,
  87, 2,
  88, 2,
  89, 2,
  90, 2,
  91, 2,
  92, 2,
  93, 2,
  94, 2,
  95, 2,
  96, 2,
  97, 2,
  98, 2,
  99, 2,
  100, 2,
  101, 2,
  102, 2,
  103, 2,
  104, 2,
  105, 2,
  106, 2,
  107, 2,
  108, 2,
  109, 2,
  110, 2,
  111, 2,
  112, 2,
  113, 2,
  114, 2,
  115, 2,
  116, 2,
  117, 2,
  118, 2,
  119, 2,
  120, 2,
  121, 2,
  122, 2,
  123, 2,
  124, 2,
  125, 2,
  126, 2,
  127, 2,
  128, 2,
  129, 2,
  130, 2,
  131, 2,
  132, 2,
  133, 2,
  134, 2,
  135, 2,
  136, 2,
  137, 2,
  138, 2,
  139, 2,
  140, 2,
  141, 2,
  142, 2,
  143, 2,
  144, 2,
  1, 3,
  2, 3,
  3, 3,
  4, 3,
  5, 3,
  6, 3,
  7, 3,
  8, 3,
  9, 3,
  10, 3,
  11, 3,
  12, 3,
  13, 3,
  14, 3,
  15, 3,
  16, 3,
  17, 3,
  18, 3,
  19, 3,
  20, 3,
  21, 3,
  22, 3,
  23, 3,
  24, 3,
  25, 3,
  26, 3,
  27, 3,
  28, 3,
  29, 3,
  30, 3,
  31, 3,
  32, 3,
  33, 3,
  34, 3,
  35, 3,
  36, 3,
  37, 3,
  38, 3,
  39, 3,
  40, 3,
  41, 3,
  42, 3,
  43, 3,
  44, 3,
  45, 3,
  46, 3,
  47, 3,
  48, 3,
  49, 3,
  50, 3,
  51, 3,
  52, 3,
  53, 3,
  54, 3,
  55, 3,
  56, 3,
  57, 3,
  58, 3,
  59, 3,
  60, 3,
  61, 3,
  62, 3,
  63, 3,
  64, 3,
  65, 3,
  66, 3,
  67, 3,
  68, 3,
  69, 3,
  70, 3,
  71, 3,
  72, 3,
  73, 3,
  74, 3,
  75, 3,
  76, 3,
  77, 3,
  78, 3,
  79, 3,
  80, 3,
  81, 3,
  82, 3,
  83, 3,
  84, 3,
  85, 3,
  86, 3,
  87, 3,
  88, 3,
  89, 3,
  90, 3,
  91, 3,
  92, 3,
  93, 3,
  94, 3,
  95, 3,
  96, 3,
  97, 3,
  98, 3,
  99, 3,
  100, 3,
  101, 3,
  102, 3,
  103, 3,
  104, 3,
  105, 3,
  106, 3,
  107, 3,
  108, 3,
  109, 3,
  110, 3,
  111, 3,
  112, 3,
  113, 3,
  114, 3,
  115, 3,
  116, 3,
  117, 3,
  118, 3,
  119, 3,
  120, 3,
  121, 3,
  122, 3,
  123, 3,
  124, 3,
  125, 3,
  126, 3,
  127, 3,
  128, 3,
  129, 3,
  130, 3,
  131, 3,
  132, 3,
  133, 3,
  134, 3,
  135, 3,
  136, 3,
  137, 3,
  138, 3,
  139, 3,
  140, 3,
  141, 3,
  142, 3,
  143, 3,
  144, 3,
  1, 4,
  2, 4,
  3, 4,
  4, 4,
  5, 4,
  6, 4,
  7, 4,
  8, 4,
  9, 4,
  10, 4,
  11, 4,
  12, 4,
  13, 4,
  14, 4,
  15, 4,
  16, 4,
  17, 4,
  18, 4,
  19, 4,
  20, 4,
  21, 4,
  22, 4,
  23, 4,
  24, 4,
  25, 4,
  26, 4,
  27, 4,
  28, 4,
  29, 4,
  30, 4,
  31, 4,
  32, 4,
  33, 4,
  34, 4,
  35, 4,
  36, 4,
  37, 4,
  38, 4,
  39, 4,
  40, 4,
  41, 4,
  42, 4,
  43, 4,
  44, 4,
  45, 4,
  46, 4,
  47, 4,
  48, 4,
  49, 4,
  50, 4,
  51, 4,
  52, 4,
  53, 4,
  54, 4,
  55, 4,
  56, 4,
  57, 4,
  58, 4,
  59, 4,
  60, 4,
  61, 4,
  62, 4,
  63, 4,
  64, 4,
  65, 4,
  66, 4,
  67, 4,
  68, 4,
  69, 4,
  70, 4,
  71, 4,
  72, 4,
  73, 4,
  74, 4,
  75, 4,
  76, 4,
  77, 4,
  78, 4,
  79, 4,
  80, 4,
  81, 4,
  82, 4,
  83, 4,
  84, 4,
  85, 4,
  86, 4,
  87, 4,
  88, 4,
  89, 4,
  90, 4,
  91, 4,
  92, 4,
  93, 4,
  94, 4,
  95, 4,
  96, 4,
  97, 4,
  98, 4,
  99, 4,
  100, 4,
  101, 4,
  102, 4,
  103, 4,
  104, 4,
  105, 4,
  106, 4,
  107, 4,
  108, 4,
  109, 4,
  110, 4,
  111, 4,
  112, 4,
  113, 4,
  114, 4,
  115, 4,
  116, 4,
  117, 4,
  118, 4,
  119, 4,
  120, 4,
  121, 4,
  122, 4,
  123, 4,
  124, 4,
  125, 4,
  126, 4,
  127, 4,
  128, 4,
  129, 4,
  130, 4,
  131, 4,
  132, 4,
  133, 4,
  134, 4,
  135, 4,
  136, 4,
  137, 4,
  138, 4,
  139, 4,
  140, 4,
  141, 4,
  142, 4,
  143, 4,
  144, 4,
  1, 5,
  2, 5,
  3, 5,
  4, 5,
  5, 5,
  6, 5,
  7, 5,
  8, 5,
  9, 5,
  10, 5,
  11, 5,
  12, 5,
  13, 5,
  14, 5,
  15, 5,
  16, 5,
  17, 5,
  18, 5,
  19, 5,
  20, 5,
  21, 5,
  22, 5,
  23, 5,
  24, 5,
  25, 5,
  26, 5,
  27, 5,
  28, 5,
  29, 5,
  30, 5,
  31, 5,
  32, 5,
  33, 5,
  34, 5,
  35, 5,
  36, 5,
  37, 5,
  38, 5,
  39, 5,
  40, 5,
  41, 5,
  42, 5,
  43, 5,
  44, 5,
  45, 5,
  46, 5,
  47, 5,
  48, 5,
  49, 5,
  50, 5,
  51, 5,
  52, 5,
  53, 5,
  54, 5,
  55, 5,
  56, 5,
  57, 5,
  58, 5,
  59, 5,
  60, 5,
  61, 5,
  62, 5,
  63, 5,
  64, 5,
  65, 5,
  66, 5,
  67, 5,
  68, 5,
  69, 5,
  70, 5,
  71, 5,
  72, 5,
  73, 5,
  74, 5,
  75, 5,
  76, 5,
  77, 5,
  78, 5,
  79, 5,
  80, 5,
  81, 5,
  82, 5,
  83, 5,
  84, 5,
  85, 5,
  86, 5,
  87, 5,
  88, 5,
  89, 5,
  90, 5,
  91, 5,
  92, 5,
  93, 5,
  94, 5,
  95, 5,
  96, 5,
  97, 5,
  98, 5,
  99, 5,
  100, 5,
  101, 5,
  102, 5,
  103, 5,
  104, 5,
  105, 5,
  106, 5,
  107, 5,
  108, 5,
  109, 5,
  110, 5,
  111, 5,
  112, 5,
  113, 5,
  114, 5,
  115, 5,
  116, 5,
  117, 5,
  118, 5,
  119, 5,
  120, 5,
  121, 5,
  122, 5,
  123, 5,
  124, 5,
  125, 5,
  126, 5,
  127, 5,
  128, 5,
  129, 5,
  130, 5,
  131, 5,
  132, 5,
  133, 5,
  134, 5,
  135, 5,
  136, 5,
  137, 5,
  138, 5,
  139, 5,
  140, 5,
  141, 5,
  142, 5,
  143, 5,
  144, 5,
  1, 6,
  2, 6,
  3, 6,
  4, 6,
  5, 6,
  6, 6,
  7, 6,
  8, 6,
  9, 6,
  10, 6,
  11, 6,
  12, 6,
  13, 6,
  14, 6,
  15, 6,
  16, 6,
  17, 6,
  18, 6,
  19, 6,
  20, 6,
  21, 6,
  22, 6,
  23, 6,
  24, 6,
  25, 6,
  26, 6,
  27, 6,
  28, 6,
  29, 6,
  30, 6,
  31, 6,
  32, 6,
  33, 6,
  34, 6,
  35, 6,
  36, 6,
  37, 6,
  38, 6,
  39, 6,
  40, 6,
  41, 6,
  42, 6,
  43, 6,
  44, 6,
  45, 6,
  46, 6,
  47, 6,
  48, 6,
  49, 6,
  50, 6,
  51, 6,
  52, 6,
  53, 6,
  54, 6,
  55, 6,
  56, 6,
  57, 6,
  58, 6,
  59, 6,
  60, 6,
  61, 6,
  62, 6,
  63, 6,
  64, 6,
  65, 6,
  66, 6,
  67, 6,
  68, 6,
  69, 6,
  70, 6,
  71, 6,
  72, 6,
  73, 6,
  74, 6,
  75, 6,
  76, 6,
  77, 6,
  78, 6,
  79, 6,
  80, 6,
  81, 6,
  82, 6,
  83, 6,
  84, 6,
  85, 6,
  86, 6,
  87, 6,
  88, 6,
  89, 6,
  90, 6,
  91, 6,
  92, 6,
  93, 6,
  94, 6,
  95, 6,
  96, 6,
  97, 6,
  98, 6,
  99, 6,
  100, 6,
  101, 6,
  102, 6,
  103, 6,
  104, 6,
  105, 6,
  106, 6,
  107, 6,
  108, 6,
  109, 6,
  110, 6,
  111, 6,
  112, 6,
  113, 6,
  114, 6,
  115, 6,
  116, 6,
  117, 6,
  118, 6,
  119, 6,
  120, 6,
  121, 6,
  122, 6,
  123, 6,
  124, 6,
  125, 6,
  126, 6,
  127, 6,
  128, 6,
  129, 6,
  130, 6,
  131, 6,
  132, 6,
  133, 6,
  134, 6,
  135, 6,
  136, 6,
  137, 6,
  138, 6,
  139, 6,
  140, 6,
  141, 6,
  142, 6,
  143, 6,
  144, 6,
  1, 7,
  2, 7,
  3, 7,
  4, 7,
  5, 7,
  6, 7,
  7, 7,
  8, 7,
  9, 7,
  10, 7,
  11, 7,
  12, 7,
  13, 7,
  14, 7,
  15, 7,
  16, 7,
  17, 7,
  18, 7,
  19, 7,
  20, 7,
  21, 7,
  22, 7,
  23, 7,
  24, 7,
  25, 7,
  26, 7,
  27, 7,
  28, 7,
  29, 7,
  30, 7,
  31, 7,
  32, 7,
  33, 7,
  34, 7,
  35, 7,
  36, 7,
  37, 7,
  38, 7,
  39, 7,
  40, 7,
  41, 7,
  42, 7,
  43, 7,
  44, 7,
  45, 7,
  46, 7,
  47, 7,
  48, 7,
  49, 7,
  50, 7,
  51, 7,
  52, 7,
  53, 7,
  54, 7,
  55, 7,
  56, 7,
  57, 7,
  58, 7,
  59, 7,
  60, 7,
  61, 7,
  62, 7,
  63, 7,
  64, 7,
  65, 7,
  66, 7,
  67, 7,
  68, 7,
  69, 7,
  70, 7,
  71, 7,
  72, 7,
  73, 7,
  74, 7,
  75, 7,
  76, 7,
  77, 7,
  78, 7,
  79, 7,
  80, 7,
  81, 7,
  82, 7,
  83, 7,
  84, 7,
  85, 7,
  86, 7,
  87, 7,
  88, 7,
  89, 7,
  90, 7,
  91, 7,
  92, 7,
  93, 7,
  94, 7,
  95, 7,
  96, 7,
  97, 7,
  98, 7,
  99, 7,
  100, 7,
  101, 7,
  102, 7,
  103, 7,
  104, 7,
  105, 7,
  106, 7,
  107, 7,
  108, 7,
  109, 7,
  110, 7,
  111, 7,
  112, 7,
  113, 7,
  114, 7,
  115, 7,
  116, 7,
  117, 7,
  118, 7,
  119, 7,
  120, 7,
  121, 7,
  122, 7,
  123, 7,
  124, 7,
  125, 7,
  126, 7,
  127, 7,
  128, 7,
  129, 7,
  130, 7,
  131, 7,
  132, 7,
  133, 7,
  134, 7,
  135, 7,
  136, 7,
  137, 7,
  138, 7,
  139, 7,
  140, 7,
  141, 7,
  142, 7,
  143, 7,
  144, 7,
  1, 8,
  2, 8,
  3, 8,
  4, 8,
  5, 8,
  6, 8,
  7, 8,
  8, 8,
  9, 8,
  10, 8,
  11, 8,
  12, 8,
  13, 8,
  14, 8,
  15, 8,
  16, 8,
  17, 8,
  18, 8,
  19, 8,
  20, 8,
  21, 8,
  22, 8,
  23, 8,
  24, 8,
  25, 8,
  26, 8,
  27, 8,
  28, 8,
  29, 8,
  30, 8,
  31, 8,
  32, 8,
  33, 8,
  34, 8,
  35, 8,
  36, 8,
  37, 8,
  38, 8,
  39, 8,
  40, 8,
  41, 8,
  42, 8,
  43, 8,
  44, 8,
  45, 8,
  46, 8,
  47, 8,
  48, 8,
  49, 8,
  50, 8,
  51, 8,
  52, 8,
  53, 8,
  54, 8,
  55, 8,
  56, 8,
  57, 8,
  58, 8,
  59, 8,
  60, 8,
  61, 8,
  62, 8,
  63, 8,
  64, 8,
  65, 8,
  66, 8,
  85, 8,
  86, 8,
  87, 8,
  88, 8,
  89, 8,
  90, 8,
  91, 8,
  92, 8,
  93, 8,
  94, 8,
  95, 8,
  96, 8,
  97, 8,
  98, 8,
  99, 8,
  100, 8,
  101, 8,
  102, 8,
  103, 8,
  104, 8,
  105, 8,
  106, 8,
  107, 8,
  108, 8,
  109, 8,
  110, 8,
  111, 8,
  112, 8,
  113, 8,
  114, 8,
  115, 8,
  116, 8,
  117, 8,
  118, 8,
  119, 8,
  120, 8,
  121, 8,
  122, 8,
  123, 8,
  133, 8,
  134, 8,
  135, 8,
  136, 8,
  137, 8,
  138, 8,
  139, 8,
  140, 8,
  141, 8,
  142, 8,
  143, 8,
  144, 8,
  1, 9,
  2, 9,
  3, 9,
  4, 9,
  5, 9,
  6, 9,
  7, 9,
  8, 9,
  9, 9,
  10, 9,
  11, 9,
  12, 9,
  13, 9,
  14, 9,
  15, 9,
  16, 9,
  17, 9,
  18, 9,
  19, 9,
  20, 9,
  21, 9,
  22, 9,
  23, 9,
  24, 9,
  25, 9,
  26, 9,
  27, 9,
  28, 9,
  29, 9,
  30, 9,
  31, 9,
  32, 9,
  33, 9,
  34, 9,
  35, 9,
  36, 9,
  37, 9,
  38, 9,
  39, 9,
  40, 9,
  41, 9,
  42, 9,
  43, 9,
  44, 9,
  45, 9,
  46, 9,
  47, 9,
  48, 9,
  49, 9,
  50, 9,
  51, 9,
  52, 9,
  53, 9,
  54, 9,
  55, 9,
  56, 9,
  57, 9,
  58, 9,
  59, 9,
  60, 9,
  61, 9,
  62, 9,
  63, 9,
  64, 9,
  65, 9,
  66, 9,
  67, 9,
  68, 9,
  91, 9,
  92, 9,
  93, 9,
  94, 9,
  95, 9,
  96, 9,
  97, 9,
  98, 9,
  99, 9,
  100, 9,
  101, 9,
  102, 9,
  103, 9,
  104, 9,
  105, 9,
  106, 9,
  107, 9,
  108, 9,
  109, 9,
  110, 9,
  111, 9,
  112, 9,
  113, 9,
  114, 9,
  115, 9,
  116, 9,
  117, 9,
  118, 9,
  119, 9,
  120, 9,
  121, 9,
  136, 9,
  137, 9,
  138, 9,
  139, 9,
  140, 9,
  141, 9,
  142, 9,
  143, 9,
  144, 9,
  1, 10,
  2, 10,
  3, 10,
  4, 10,
  5, 10,
  6, 10,
  7, 10,
  8, 10,
  9, 10,
  10, 10,
  11, 10,
  12, 10,
  13, 10,
  14, 10,
  15, 10,
  16, 10,
  17, 10,
  18, 10,
  19, 10,
  20, 10,
  21, 10,
  22, 10,
  23, 10,
  24, 10,
  25, 10,
  26, 10,
  27, 10,
  28, 10,
  29, 10,
  30, 10,
  31, 10,
  32, 10,
  33, 10,
  34, 10,
  35, 10,
  36, 10,
  37, 10,
  38, 10,
  39, 10,
  40, 10,
  41, 10,
  42, 10,
  43, 10,
  44, 10,
  45, 10,
  46, 10,
  47, 10,
  48, 10,
  49, 10,
  50, 10,
  51, 10,
  52, 10,
  53, 10,
  54, 10,
  55, 10,
  56, 10,
  57, 10,
  58, 10,
  59, 10,
  60, 10,
  61, 10,
  62, 10,
  63, 10,
  64, 10,
  65, 10,
  66, 10,
  67, 10,
  68, 10,
  69, 10,
  104, 10,
  105, 10,
  106, 10,
  107, 10,
  108, 10,
  113, 10,
  114, 10,
  115, 10,
  116, 10,
  117, 10,
  118, 10,
  119, 10,
  120, 10,
  138, 10,
  139, 10,
  140, 10,
  141, 10,
  142, 10,
  143, 10,
  144, 10,
  1, 11,
  2, 11,
  3, 11,
  4, 11,
  5, 11,
  6, 11,
  7, 11,
  8, 11,
  9, 11,
  10, 11,
  11, 11,
  12, 11,
  13, 11,
  14, 11,
  15, 11,
  16, 11,
  17, 11,
  18, 11,
  19, 11,
  20, 11,
  21, 11,
  22, 11,
  23, 11,
  24, 11,
  25, 11,
  26, 11,
  27, 11,
  28, 11,
  29, 11,
  30, 11,
  31, 11,
  32, 11,
  33, 11,
  34, 11,
  35, 11,
  36, 11,
  37, 11,
  38, 11,
  39, 11,
  40, 11,
  41, 11,
  42, 11,
  43, 11,
  44, 11,
  45, 11,
  46, 11,
  47, 11,
  48, 11,
  49, 11,
  50, 11,
  51, 11,
  52, 11,
  53, 11,
  54, 11,
  55, 11,
  56, 11,
  57, 11,
  58, 11,
  59, 11,
  60, 11,
  61, 11,
  62, 11,
  63, 11,
  64, 11,
  65, 11,
  66, 11,
  67, 11,
  114, 11,
  115, 11,
  116, 11,
  117, 11,
  118, 11,
  119, 11,
  120, 11,
  143, 11,
  144, 11,
  14, 12,
  17, 12,
  18, 12,
  19, 12,
  20, 12,
  21, 12,
  22, 12,
  23, 12,
  24, 12,
  25, 12,
  26, 12,
  27, 12,
  28, 12,
  32, 12,
  33, 12,
  34, 12,
  35, 12,
  36, 12,
  37, 12,
  38, 12,
  39, 12,
  40, 12,
  41, 12,
  42, 12,
  43, 12,
  44, 12,
  45, 12,
  46, 12,
  47, 12,
  48, 12,
  49, 12,
  50, 12,
  51, 12,
  52, 12,
  53, 12,
  54, 12,
  55, 12,
  56, 12,
  57, 12,
  58, 12,
  59, 12,
  60, 12,
  61, 12,
  62, 12,
  117, 12,
  118, 12,
  119, 12,
  120, 12,
  21, 13,
  22, 13,
  23, 13,
  35, 13,
  36, 13,
  38, 13,
  39, 13,
  40, 13,
  41, 13,
  42, 13,
  43, 13,
  44, 13,
  45, 13,
  46, 13,
  47, 13,
  51, 13,
  53, 13,
  54, 13,
  55, 13,
  56, 13,
  118, 13,
  119, 13,
  120, 13,
  121, 13,
  122, 13,
  119, 14,
  120, 14,
  121, 14,
  122, 14,
  115, 18,
  116, 18,
  117, 18,
  118, 18,
  115, 19,
  116, 19,
  117, 19,
  118, 19,
  114, 20,
  115, 20,
  116, 20,
  117, 20,
  120, 20,
  121, 20,
  28, 21,
  114, 21,
  115, 21,
  116, 21,
  117, 21,
  118, 21,
  68, 22,
  114, 22,
  115, 22,
  116, 22,
  117, 22,
  118, 22,
  67, 23,
  68, 23,
  69, 23,
  115, 23,
  116, 23,
  117, 23,
  118, 23,
  59, 24,
  60, 24,
  68, 24,
  69, 24,
  70, 24,
  115, 24,
  116, 24,
  117, 24,
  118, 24,
  59, 25,
  60, 25,
  69, 25,
  70, 25,
  71, 25,
  115, 25,
  116, 25,
  117, 25,
  118, 25,
  119, 25,
  120, 25,
  58, 26,
  59, 26,
  70, 26,
  71, 26,
  72, 26,
  115, 26,
  116, 26,
  117, 26,
  118, 26,
  119, 26,
  120, 26,
  121, 26,
  57, 27,
  58, 27,
  59, 27,
  60, 27,
  70, 27,
  71, 27,
  72, 27,
  115, 27,
  116, 27,
  117, 27,
  118, 27,
  119, 27,
  120, 27,
  121, 27,
  122, 27,
  47, 28,
  48, 28,
  55, 28,
  56, 28,
  57, 28,
  58, 28,
  59, 28,
  60, 28,
  61, 28,
  70, 28,
  115, 28,
  116, 28,
  117, 28,
  118, 28,
  119, 28,
  120, 28,
  121, 28,
  122, 28,
  123, 28,
  8, 29,
  9, 29,
  10, 29,
  11, 29,
  12, 29,
  47, 29,
  48, 29,
  49, 29,
  50, 29,
  51, 29,
  54, 29,
  55, 29,
  56, 29,
  57, 29,
  58, 29,
  59, 29,
  60, 29,
  61, 29,
  116, 29,
  117, 29,
  118, 29,
  119, 29,
  120, 29,
  121, 29,
  122, 29,
  123, 29,
  124, 29,
  7, 30,
  8, 30,
  9, 30,
  10, 30,
  11, 30,
  12, 30,
  13, 30,
  47, 30,
  48, 30,
  49, 30,
  50, 30,
  51, 30,
  52, 30,
  53, 30,
  54, 30,
  55, 30,
  56, 30,
  57, 30,
  58, 30,
  59, 30,
  60, 30,
  61, 30,
  62, 30,
  116, 30,
  117, 30,
  118, 30,
  119, 30,
  120, 30,
  121, 30,
  122, 30,
  123, 30,
  124, 30,
  7, 31,
  8, 31,
  9, 31,
  10, 31,
  11, 31,
  12, 31,
  13, 31,
  47, 31,
  48, 31,
  49, 31,
  50, 31,
  51, 31,
  52, 31,
  53, 31,
  54, 31,
  55, 31,
  56, 31,
  57, 31,
  58, 31,
  59, 31,
  60, 31,
  61, 31,
  62, 31,
  116, 31,
  117, 31,
  118, 31,
  119, 31,
  120, 31,
  121, 31,
  122, 31,
  123, 31,
  124, 31,
  125, 31,
  7, 32,
  8, 32,
  9, 32,
  10, 32,
  11, 32,
  12, 32,
  13, 32,
  14, 32,
  46, 32,
  47, 32,
  48, 32,
  49, 32,
  50, 32,
  51, 32,
  52, 32,
  53, 32,
  54, 32,
  55, 32,
  56, 32,
  57, 32,
  58, 32,
  59, 32,
  60, 32,
  61, 32,
  62, 32,
  116, 32,
  117, 32,
  118, 32,
  119, 32,
  120, 32,
  121, 32,
  122, 32,
  123, 32,
  124, 32,
  125, 32,
  7, 33,
  8, 33,
  9, 33,
  10, 33,
  11, 33,
  12, 33,
  13, 33,
  14, 33,
  18, 33,
  19, 33,
  46, 33,
  47, 33,
  48, 33,
  49, 33,
  50, 33,
  51, 33,
  52, 33,
  53, 33,
  54, 33,
  55, 33,
  56, 33,
  57, 33,
  58, 33,
  59, 33,
  60, 33,
  61, 33,
  62, 33,
  116, 33,
  117, 33,
  118, 33,
  119, 33,
  120, 33,
  121, 33,
  122, 33,
  123, 33,
  124, 33,
  125, 33,
  126, 33,
  6, 34,
  7, 34,
  8, 34,
  9, 34,
  10, 34,
  11, 34,
  12, 34,
  13, 34,
  14, 34,
  18, 34,
  19, 34,
  20, 34,
  46, 34,
  47, 34,
  48, 34,
  49, 34,
  50, 34,
  51, 34,
  52, 34,
  53, 34,
  54, 34,
  55, 34,
  56, 34,
  57, 34,
  58, 34,
  59, 34,
  60, 34,
  61, 34,
  116, 34,
  117, 34,
  118, 34,
  119, 34,
  120, 34,
  121, 34,
  122, 34,
  123, 34,
  124, 34,
  125, 34,
  126, 34,
  127, 34,
  128, 34,
  6, 35,
  7, 35,
  8, 35,
  9, 35,
  10, 35,
  11, 35,
  12, 35,
  13, 35,
  14, 35,
  18, 35,
  19, 35,
  20, 35,
  23, 35,
  46, 35,
  47, 35,
  48, 35,
  49, 35,
  50, 35,
  51, 35,
  52, 35,
  53, 35,
  54, 35,
  55, 35,
  56, 35,
  57, 35,
  58, 35,
  59, 35,
  60, 35,
  61, 35,
  67, 35,
  117, 35,
  118, 35,
  119, 35,
  120, 35,
  121, 35,
  122, 35,
  123, 35,
  124, 35,
  125, 35,
  126, 35,
  127, 35,
  128, 35,
  5, 36,
  6, 36,
  7, 36,
  8, 36,
  9, 36,
  10, 36,
  11, 36,
  12, 36,
  13, 36,
  14, 36,
  15, 36,
  18, 36,
  19, 36,
  20, 36,
  48, 36,
  49, 36,
  50, 36,
  51, 36,
  52, 36,
  53, 36,
  54, 36,
  55, 36,
  56, 36,
  57, 36,
  58, 36,
  59, 36,
  60, 36,
  117, 36,
  118, 36,
  119, 36,
  120, 36,
  121, 36,
  122, 36,
  123, 36,
  124, 36,
  125, 36,
  126, 36,
  127, 36,
  128, 36,
  5, 37,
  6, 37,
  7, 37,
  8, 37,
  9, 37,
  10, 37,
  11, 37,
  12, 37,
  13, 37,
  14, 37,
  15, 37,
  16, 37,
  18, 37,
  19, 37,
  20, 37,
  49, 37,
  50, 37,
  51, 37,
  52, 37,
  53, 37,
  54, 37,
  55, 37,
  56, 37,
  57, 37,
  58, 37,
  59, 37,
  71, 37,
  72, 37,
  115, 37,
  116, 37,
  117, 37,
  118, 37,
  119, 37,
  120, 37,
  121, 37,
  122, 37,
  123, 37,
  124, 37,
  125, 37,
  126, 37,
  127, 37,
  128, 37,
  129, 37,
  5, 38,
  6, 38,
  7, 38,
  8, 38,
  9, 38,
  10, 38,
  11, 38,
  12, 38,
  13, 38,
  14, 38,
  15, 38,
  16, 38,
  19, 38,
  20, 38,
  50, 38,
  51, 38,
  52, 38,
  53, 38,
  54, 38,
  55, 38,
  57, 38,
  58, 38,
  59, 38,
  114, 38,
  115, 38,
  116, 38,
  117, 38,
  118, 38,
  119, 38,
  120, 38,
  121, 38,
  122, 38,
  123, 38,
  124, 38,
  125, 38,
  126, 38,
  127, 38,
  128, 38,
  129, 38,
  5, 39,
  6, 39,
  7, 39,
  8, 39,
  9, 39,
  10, 39,
  11, 39,
  12, 39,
  13, 39,
  14, 39,
  15, 39,
  16, 39,
  20, 39,
  51, 39,
  52, 39,
  53, 39,
  54, 39,
  55, 39,
  57, 39,
  58, 39,
  114, 39,
  115, 39,
  116, 39,
  117, 39,
  118, 39,
  119, 39,
  120, 39,
  121, 39,
  122, 39,
  123, 39,
  124, 39,
  125, 39,
  126, 39,
  127, 39,
  128, 39,
  129, 39,
  6, 40,
  7, 40,
  8, 40,
  9, 40,
  10, 40,
  11, 40,
  12, 40,
  13, 40,
  14, 40,
  15, 40,
  16, 40,
  50, 40,
  53, 40,
  54, 40,
  55, 40,
  57, 40,
  58, 40,
  61, 40,
  113, 40,
  114, 40,
  115, 40,
  116, 40,
  117, 40,
  118, 40,
  119, 40,
  120, 40,
  121, 40,
  122, 40,
  123, 40,
  124, 40,
  125, 40,
  126, 40,
  127, 40,
  128, 40,
  129, 40,
  130, 40,
  6, 41,
  7, 41,
  8, 41,
  9, 41,
  10, 41,
  11, 41,
  12, 41,
  13, 41,
  14, 41,
  15, 41,
  16, 41,
  47, 41,
  48, 41,
  49, 41,
  50, 41,
  51, 41,
  57, 41,
  58, 41,
  59, 41,
  60, 41,
  61, 41,
  113, 41,
  114, 41,
  115, 41,
  116, 41,
  117, 41,
  118, 41,
  119, 41,
  120, 41,
  121, 41,
  122, 41,
  123, 41,
  124, 41,
  125, 41,
  126, 41,
  127, 41,
  128, 41,
  129, 41,
  130, 41,
  5, 42,
  6, 42,
  7, 42,
  8, 42,
  9, 42,
  10, 42,
  11, 42,
  12, 42,
  13, 42,
  14, 42,
  15, 42,
  16, 42,
  43, 42,
  44, 42,
  45, 42,
  46, 42,
  47, 42,
  48, 42,
  49, 42,
  53, 42,
  54, 42,
  56, 42,
  57, 42,
  58, 42,
  59, 42,
  60, 42,
  61, 42,
  63, 42,
  112, 42,
  113, 42,
  114, 42,
  115, 42,
  116, 42,
  117, 42,
  118, 42,
  119, 42,
  120, 42,
  121, 42,
  122, 42,
  123, 42,
  124, 42,
  125, 42,
  126, 42,
  127, 42,
  128, 42,
  129, 42,
  130, 42,
  5, 43,
  6, 43,
  7, 43,
  8, 43,
  9, 43,
  10, 43,
  11, 43,
  12, 43,
  13, 43,
  14, 43,
  15, 43,
  16, 43,
  41, 43,
  42, 43,
  43, 43,
  48, 43,
  49, 43,
  50, 43,
  54, 43,
  55, 43,
  56, 43,
  57, 43,
  58, 43,
  59, 43,
  60, 43,
  61, 43,
  112, 43,
  113, 43,
  114, 43,
  115, 43,
  116, 43,
  117, 43,
  118, 43,
  119, 43,
  120, 43,
  121, 43,
  122, 43,
  123, 43,
  124, 43,
  125, 43,
  126, 43,
  127, 43,
  128, 43,
  129, 43,
  130, 43,
  4, 44,
  5, 44,
  6, 44,
  7, 44,
  8, 44,
  9, 44,
  10, 44,
  11, 44,
  12, 44,
  13, 44,
  14, 44,
  15, 44,
  16, 44,
  17, 44,
  41, 44,
  42, 44,
  43, 44,
  45, 44,
  46, 44,
  47, 44,
  48, 44,
  49, 44,
  50, 44,
  51, 44,
  52, 44,
  53, 44,
  54, 44,
  55, 44,
  56, 44,
  57, 44,
  58, 44,
  112, 44,
  113, 44,
  114, 44,
  115, 44,
  116, 44,
  117, 44,
  118, 44,
  119, 44,
  120, 44,
  121, 44,
  122, 44,
  123, 44,
  124, 44,
  125, 44,
  126, 44,
  127, 44,
  128, 44,
  129, 44,
  4, 45,
  5, 45,
  6, 45,
  7, 45,
  8, 45,
  9, 45,
  10, 45,
  11, 45,
  12, 45,
  13, 45,
  14, 45,
  15, 45,
  16, 45,
  17, 45,
  18, 45,
  41, 45,
  42, 45,
  43, 45,
  44, 45,
  45, 45,
  46, 45,
  47, 45,
  48, 45,
  49, 45,
  50, 45,
  51, 45,
  52, 45,
  53, 45,
  54, 45,
  55, 45,
  56, 45,
  112, 45,
  113, 45,
  114, 45,
  115, 45,
  116, 45,
  117, 45,
  118, 45,
  119, 45,
  120, 45,
  121, 45,
  122, 45,
  123, 45,
  124, 45,
  125, 45,
  126, 45,
  4, 46,
  5, 46,
  6, 46,
  7, 46,
  8, 46,
  9, 46,
  10, 46,
  11, 46,
  12, 46,
  13, 46,
  14, 46,
  15, 46,
  16, 46,
  17, 46,
  18, 46,
  39, 46,
  40, 46,
  41, 46,
  42, 46,
  44, 46,
  45, 46,
  46, 46,
  47, 46,
  48, 46,
  49, 46,
  50, 46,
  51, 46,
  52, 46,
  113, 46,
  114, 46,
  115, 46,
  116, 46,
  117, 46,
  118, 46,
  119, 46,
  120, 46,
  121, 46,
  122, 46,
  123, 46,
  124, 46,
  4, 47,
  5, 47,
  6, 47,
  7, 47,
  8, 47,
  9, 47,
  10, 47,
  11, 47,
  12, 47,
  13, 47,
  14, 47,
  15, 47,
  16, 47,
  17, 47,
  18, 47,
  19, 47,
  20, 47,
  39, 47,
  40, 47,
  41, 47,
  42, 47,
  44, 47,
  45, 47,
  46, 47,
  47, 47,
  48, 47,
  52, 47,
  113, 47,
  114, 47,
  115, 47,
  116, 47,
  117, 47,
  118, 47,
  119, 47,
  120, 47,
  121, 47,
  122, 47,
  123, 47,
  124, 47,
  1, 48,
  3, 48,
  4, 48,
  5, 48,
  6, 48,
  7, 48,
  8, 48,
  9, 48,
  10, 48,
  11, 48,
  12, 48,
  13, 48,
  14, 48,
  15, 48,
  16, 48,
  17, 48,
  18, 48,
  19, 48,
  20, 48,
  39, 48,
  40, 48,
  41, 48,
  42, 48,
  46, 48,
  47, 48,
  48, 48,
  51, 48,
  114, 48,
  115, 48,
  116, 48,
  117, 48,
  118, 48,
  119, 48,
  120, 48,
  121, 48,
  122, 48,
  123, 48,
  124, 48,
  141, 48,
  142, 48,
  143, 48,
  144, 48,
  1, 49,
  2, 49,
  3, 49,
  4, 49,
  5, 49,
  6, 49,
  7, 49,
  8, 49,
  9, 49,
  10, 49,
  11, 49,
  12, 49,
  13, 49,
  14, 49,
  15, 49,
  16, 49,
  17, 49,
  18, 49,
  19, 49,
  20, 49,
  31, 49,
  32, 49,
  33, 49,
  40, 49,
  41, 49,
  42, 49,
  47, 49,
  48, 49,
  49, 49,
  50, 49,
  51, 49,
  111, 49,
  112, 49,
  113, 49,
  114, 49,
  115, 49,
  116, 49,
  117, 49,
  118, 49,
  119, 49,
  120, 49,
  121, 49,
  122, 49,
  139, 49,
  140, 49,
  141, 49,
  142, 49,
  143, 49,
  144, 49,
  1, 50,
  2, 50,
  3, 50,
  4, 50,
  5, 50,
  6, 50,
  7, 50,
  8, 50,
  9, 50,
  10, 50,
  11, 50,
  12, 50,
  13, 50,
  14, 50,
  15, 50,
  16, 50,
  17, 50,
  18, 50,
  19, 50,
  20, 50,
  21, 50,
  31, 50,
  32, 50,
  33, 50,
  40, 50,
  42, 50,
  43, 50,
  44, 50,
  47, 50,
  48, 50,
  50, 50,
  51, 50,
  110, 50,
  111, 50,
  112, 50,
  113, 50,
  114, 50,
  115, 50,
  116, 50,
  117, 50,
  118, 50,
  119, 50,
  120, 50,
  139, 50,
  140, 50,
  141, 50,
  142, 50,
  143, 50,
  144, 50,
  1, 51,
  2, 51,
  3, 51,
  4, 51,
  5, 51,
  6, 51,
  7, 51,
  8, 51,
  9, 51,
  10, 51,
  11, 51,
  12, 51,
  13, 51,
  14, 51,
  15, 51,
  16, 51,
  17, 51,
  18, 51,
  19, 51,
  20, 51,
  21, 51,
  31, 51,
  32, 51,
  40, 51,
  41, 51,
  42, 51,
  43, 51,
  44, 51,
  48, 51,
  49, 51,
  50, 51,
  110, 51,
  111, 51,
  115, 51,
  116, 51,
  117, 51,
  118, 51,
  119, 51,
  120, 51,
  138, 51,
  139, 51,
  140, 51,
  141, 51,
  142, 51,
  143, 51,
  144, 51,
  1, 52,
  2, 52,
  3, 52,
  4, 52,
  5, 52,
  6, 52,
  7, 52,
  8, 52,
  9, 52,
  10, 52,
  11, 52,
  12, 52,
  13, 52,
  14, 52,
  15, 52,
  16, 52,
  17, 52,
  18, 52,
  19, 52,
  20, 52,
  30, 52,
  31, 52,
  32, 52,
  40, 52,
  41, 52,
  42, 52,
  43, 52,
  44, 52,
  49, 52,
  50, 52,
  108, 52,
  109, 52,
  110, 52,
  111, 52,
  138, 52,
  139, 52,
  140, 52,
  141, 52,
  142, 52,
  143, 52,
  144, 52,
  1, 53,
  2, 53,
  3, 53,
  4, 53,
  5, 53,
  6, 53,
  7, 53,
  8, 53,
  9, 53,
  10, 53,
  11, 53,
  12, 53,
  13, 53,
  14, 53,
  15, 53,
  16, 53,
  17, 53,
  18, 53,
  19, 53,
  20, 53,
  21, 53,
  30, 53,
  31, 53,
  32, 53,
  33, 53,
  40, 53,
  41, 53,
  42, 53,
  43, 53,
  44, 53,
  49, 53,
  105, 53,
  106, 53,
  107, 53,
  108, 53,
  109, 53,
  110, 53,
  111, 53,
  138, 53,
  139, 53,
  140, 53,
  141, 53,
  142, 53,
  143, 53,
  144, 53,
  1, 54,
  2, 54,
  3, 54,
  4, 54,
  5, 54,
  6, 54,
  7, 54,
  8, 54,
  9, 54,
  10, 54,
  11, 54,
  12, 54,
  13, 54,
  14, 54,
  15, 54,
  16, 54,
  17, 54,
  18, 54,
  19, 54,
  20, 54,
  21, 54,
  22, 54,
  23, 54,
  30, 54,
  31, 54,
  32, 54,
  33, 54,
  34, 54,
  38, 54,
  39, 54,
  40, 54,
  41, 54,
  42, 54,
  43, 54,
  44, 54,
  49, 54,
  103, 54,
  104, 54,
  105, 54,
  106, 54,
  107, 54,
  108, 54,
  109, 54,
  115, 54,
  116, 54,
  118, 54,
  138, 54,
  139, 54,
  140, 54,
  141, 54,
  142, 54,
  143, 54,
  144, 54,
  1, 55,
  2, 55,
  3, 55,
  4, 55,
  5, 55,
  6, 55,
  7, 55,
  8, 55,
  9, 55,
  10, 55,
  11, 55,
  12, 55,
  13, 55,
  14, 55,
  15, 55,
  16, 55,
  17, 55,
  18, 55,
  19, 55,
  20, 55,
  21, 55,
  22, 55,
  23, 55,
  24, 55,
  30, 55,
  31, 55,
  32, 55,
  33, 55,
  34, 55,
  35, 55,
  38, 55,
  39, 55,
  40, 55,
  41, 55,
  42, 55,
  43, 55,
  44, 55,
  45, 55,
  82, 55,
  103, 55,
  104, 55,
  105, 55,
  106, 55,
  108, 55,
  109, 55,
  114, 55,
  115, 55,
  116, 55,
  117, 55,
  118, 55,
  138, 55,
  139, 55,
  140, 55,
  141, 55,
  142, 55,
  143, 55,
  144, 55,
  1, 56,
  2, 56,
  3, 56,
  4, 56,
  5, 56,
  6, 56,
  7, 56,
  8, 56,
  9, 56,
  10, 56,
  11, 56,
  12, 56,
  13, 56,
  14, 56,
  15, 56,
  16, 56,
  17, 56,
  18, 56,
  19, 56,
  20, 56,
  21, 56,
  22, 56,
  23, 56,
  24, 56,
  28, 56,
  29, 56,
  30, 56,
  31, 56,
  32, 56,
  33, 56,
  34, 56,
  35, 56,
  36, 56,
  37, 56,
  38, 56,
  39, 56,
  40, 56,
  41, 56,
  42, 56,
  43, 56,
  44, 56,
  45, 56,
  46, 56,
  49, 56,
  82, 56,
  102, 56,
  103, 56,
  104, 56,
  105, 56,
  106, 56,
  109, 56,
  111, 56,
  112, 56,
  113, 56,
  114, 56,
  138, 56,
  139, 56,
  140, 56,
  141, 56,
  142, 56,
  143, 56,
  144, 56,
  1, 57,
  2, 57,
  3, 57,
  4, 57,
  5, 57,
  6, 57,
  7, 57,
  8, 57,
  9, 57,
  10, 57,
  11, 57,
  12, 57,
  13, 57,
  14, 57,
  15, 57,
  16, 57,
  17, 57,
  18, 57,
  19, 57,
  20, 57,
  21, 57,
  22, 57,
  23, 57,
  24, 57,
  27, 57,
  28, 57,
  29, 57,
  30, 57,
  31, 57,
  32, 57,
  33, 57,
  34, 57,
  35, 57,
  36, 57,
  37, 57,
  38, 57,
  39, 57,
  40, 57,
  41, 57,
  42, 57,
  43, 57,
  44, 57,
  45, 57,
  46, 57,
  47, 57,
  48, 57,
  49, 57,
  100, 57,
  101, 57,
  102, 57,
  103, 57,
  104, 57,
  105, 57,
  111, 57,
  112, 57,
  113, 57,
  138, 57,
  139, 57,
  140, 57,
  141, 57,
  142, 57,
  143, 57,
  144, 57,
  1, 58,
  2, 58,
  3, 58,
  4, 58,
  5, 58,
  6, 58,
  7, 58,
  8, 58,
  9, 58,
  10, 58,
  11, 58,
  12, 58,
  13, 58,
  14, 58,
  15, 58,
  16, 58,
  17, 58,
  18, 58,
  19, 58,
  20, 58,
  21, 58,
  22, 58,
  23, 58,
  24, 58,
  25, 58,
  26, 58,
  27, 58,
  28, 58,
  29, 58,
  30, 58,
  31, 58,
  32, 58,
  33, 58,
  34, 58,
  35, 58,
  36, 58,
  37, 58,
  38, 58,
  39, 58,
  40, 58,
  41, 58,
  42, 58,
  43, 58,
  44, 58,
  45, 58,
  46, 58,
  47, 58,
  48, 58,
  49, 58,
  99, 58,
  100, 58,
  101, 58,
  102, 58,
  103, 58,
  104, 58,
  105, 58,
  106, 58,
  112, 58,
  139, 58,
  140, 58,
  141, 58,
  142, 58,
  143, 58,
  144, 58,
  1, 59,
  2, 59,
  3, 59,
  4, 59,
  5, 59,
  6, 59,
  7, 59,
  8, 59,
  9, 59,
  10, 59,
  11, 59,
  12, 59,
  13, 59,
  14, 59,
  15, 59,
  16, 59,
  17, 59,
  18, 59,
  19, 59,
  20, 59,
  21, 59,
  22, 59,
  23, 59,
  24, 59,
  25, 59,
  26, 59,
  27, 59,
  28, 59,
  29, 59,
  30, 59,
  31, 59,
  32, 59,
  33, 59,
  34, 59,
  35, 59,
  36, 59,
  37, 59,
  38, 59,
  39, 59,
  40, 59,
  41, 59,
  42, 59,
  43, 59,
  44, 59,
  45, 59,
  46, 59,
  47, 59,
  48, 59,
  49, 59,
  99, 59,
  100, 59,
  101, 59,
  102, 59,
  103, 59,
  104, 59,
  105, 59,
  106, 59,
  111, 59,
  112, 59,
  139, 59,
  140, 59,
  141, 59,
  142, 59,
  143, 59,
  144, 59,
  1, 60,
  2, 60,
  3, 60,
  4, 60,
  5, 60,
  6, 60,
  7, 60,
  8, 60,
  9, 60,
  10, 60,
  11, 60,
  12, 60,
  13, 60,
  14, 60,
  15, 60,
  16, 60,
  17, 60,
  18, 60,
  19, 60,
  20, 60,
  21, 60,
  22, 60,
  23, 60,
  24, 60,
  25, 60,
  26, 60,
  27, 60,
  28, 60,
  29, 60,
  30, 60,
  31, 60,
  32, 60,
  33, 60,
  34, 60,
  35, 60,
  36, 60,
  37, 60,
  38, 60,
  39, 60,
  40, 60,
  41, 60,
  42, 60,
  43, 60,
  44, 60,
  45, 60,
  46, 60,
  47, 60,
  48, 60,
  49, 60,
  98, 60,
  99, 60,
  100, 60,
  101, 60,
  102, 60,
  103, 60,
  104, 60,
  105, 60,
  106, 60,
  107, 60,
  108, 60,
  109, 60,
  110, 60,
  111, 60,
  112, 60,
  140, 60,
  141, 60,
  142, 60,
  143, 60,
  144, 60,
  1, 61,
  2, 61,
  3, 61,
  4, 61,
  5, 61,
  6, 61,
  7, 61,
  8, 61,
  9, 61,
  10, 61,
  11, 61,
  12, 61,
  13, 61,
  14, 61,
  15, 61,
  16, 61,
  17, 61,
  18, 61,
  19, 61,
  20, 61,
  21, 61,
  22, 61,
  23, 61,
  24, 61,
  25, 61,
  26, 61,
  27, 61,
  28, 61,
  29, 61,
  30, 61,
  31, 61,
  32, 61,
  33, 61,
  34, 61,
  35, 61,
  36, 61,
  37, 61,
  38, 61,
  39, 61,
  40, 61,
  41, 61,
  42, 61,
  43, 61,
  44, 61,
  45, 61,
  46, 61,
  47, 61,
  48, 61,
  49, 61,
  53, 61,
  98, 61,
  99, 61,
  100, 61,
  101, 61,
  102, 61,
  103, 61,
  104, 61,
  105, 61,
  106, 61,
  107, 61,
  108, 61,
  109, 61,
  110, 61,
  111, 61,
  112, 61,
  141, 61,
  142, 61,
  143, 61,
  144, 61,
  1, 62,
  2, 62,
  3, 62,
  4, 62,
  5, 62,
  6, 62,
  9, 62,
  10, 62,
  15, 62,
  16, 62,
  17, 62,
  18, 62,
  19, 62,
  20, 62,
  21, 62,
  22, 62,
  23, 62,
  24, 62,
  25, 62,
  26, 62,
  27, 62,
  28, 62,
  29, 62,
  30, 62,
  31, 62,
  32, 62,
  33, 62,
  34, 62,
  35, 62,
  36, 62,
  37, 62,
  38, 62,
  39, 62,
  40, 62,
  41, 62,
  42, 62,
  43, 62,
  44, 62,
  45, 62,
  46, 62,
  47, 62,
  48, 62,
  49, 62,
  51, 62,
  53, 62,
  54, 62,
  55, 62,
  97, 62,
  98, 62,
  99, 62,
  100, 62,
  101, 62,
  102, 62,
  103, 62,
  104, 62,
  105, 62,
  106, 62,
  107, 62,
  108, 62,
  109, 62,
  110, 62,
  111, 62,
  112, 62,
  113, 62,
  114, 62,
  141, 62,
  142, 62,
  143, 62,
  144, 62,
  1, 63,
  2, 63,
  3, 63,
  4, 63,
  5, 63,
  12, 63,
  13, 63,
  14, 63,
  15, 63,
  16, 63,
  17, 63,
  18, 63,
  19, 63,
  20, 63,
  21, 63,
  22, 63,
  23, 63,
  24, 63,
  25, 63,
  26, 63,
  27, 63,
  28, 63,
  29, 63,
  30, 63,
  31, 63,
  32, 63,
  33, 63,
  34, 63,
  35, 63,
  36, 63,
  37, 63,
  38, 63,
  39, 63,
  40, 63,
  41, 63,
  42, 63,
  43, 63,
  44, 63,
  45, 63,
  46, 63,
  47, 63,
  48, 63,
  49, 63,
  51, 63,
  52, 63,
  53, 63,
  54, 63,
  55, 63,
  56, 63,
  57, 63,
  96, 63,
  97, 63,
  98, 63,
  99, 63,
  100, 63,
  101, 63,
  102, 63,
  103, 63,
  104, 63,
  105, 63,
  106, 63,
  107, 63,
  108, 63,
  109, 63,
  110, 63,
  111, 63,
  112, 63,
  113, 63,
  114, 63,
  142, 63,
  143, 63,
  144, 63,
  1, 64,
  2, 64,
  3, 64,
  4, 64,
  5, 64,
  6, 64,
  7, 64,
  9, 64,
  10, 64,
  11, 64,
  12, 64,
  13, 64,
  14, 64,
  15, 64,
  16, 64,
  17, 64,
  18, 64,
  19, 64,
  20, 64,
  21, 64,
  22, 64,
  23, 64,
  24, 64,
  25, 64,
  26, 64,
  27, 64,
  28, 64,
  29, 64,
  30, 64,
  31, 64,
  32, 64,
  33, 64,
  34, 64,
  35, 64,
  36, 64,
  37, 64,
  38, 64,
  39, 64,
  40, 64,
  41, 64,
  42, 64,
  43, 64,
  44, 64,
  45, 64,
  46, 64,
  47, 64,
  48, 64,
  49, 64,
  51, 64,
  52, 64,
  55, 64,
  56, 64,
  57, 64,
  95, 64,
  96, 64,
  97, 64,
  98, 64,
  99, 64,
  100, 64,
  101, 64,
  102, 64,
  103, 64,
  104, 64,
  105, 64,
  106, 64,
  107, 64,
  108, 64,
  109, 64,
  110, 64,
  111, 64,
  112, 64,
  113, 64,
  114, 64,
  141, 64,
  142, 64,
  143, 64,
  144, 64,
  1, 65,
  4, 65,
  6, 65,
  7, 65,
  8, 65,
  9, 65,
  10, 65,
  11, 65,
  12, 65,
  13, 65,
  14, 65,
  15, 65,
  16, 65,
  17, 65,
  18, 65,
  19, 65,
  20, 65,
  21, 65,
  22, 65,
  23, 65,
  24, 65,
  25, 65,
  26, 65,
  27, 65,
  28, 65,
  29, 65,
  30, 65,
  31, 65,
  32, 65,
  33, 65,
  34, 65,
  35, 65,
  36, 65,
  37, 65,
  38, 65,
  39, 65,
  40, 65,
  41, 65,
  42, 65,
  43, 65,
  44, 65,
  45, 65,
  46, 65,
  47, 65,
  48, 65,
  49, 65,
  50, 65,
  51, 65,
  52, 65,
  56, 65,
  57, 65,
  95, 65,
  96, 65,
  97, 65,
  98, 65,
  99, 65,
  100, 65,
  101, 65,
  102, 65,
  103, 65,
  104, 65,
  105, 65,
  106, 65,
  107, 65,
  108, 65,
  109, 65,
  110, 65,
  111, 65,
  112, 65,
  113, 65,
  114, 65,
  115, 65,
  141, 65,
  142, 65,
  143, 65,
  144, 65,
  1, 66,
  2, 66,
  4, 66,
  5, 66,
  6, 66,
  7, 66,
  8, 66,
  9, 66,
  10, 66,
  11, 66,
  12, 66,
  13, 66,
  14, 66,
  15, 66,
  16, 66,
  17, 66,
  18, 66,
  19, 66,
  20, 66,
  21, 66,
  22, 66,
  23, 66,
  24, 66,
  25, 66,
  26, 66,
  27, 66,
  28, 66,
  29, 66,
  30, 66,
  31, 66,
  32, 66,
  33, 66,
  34, 66,
  35, 66,
  36, 66,
  37, 66,
  38, 66,
  39, 66,
  40, 66,
  41, 66,
  42, 66,
  43, 66,
  44, 66,
  45, 66,
  46, 66,
  47, 66,
  48, 66,
  49, 66,
  50, 66,
  51, 66,
  52, 66,
  53, 66,
  57, 66,
  58, 66,
  95, 66,
  96, 66,
  97, 66,
  98, 66,
  99, 66,
  100, 66,
  101, 66,
  102, 66,
  103, 66,
  104, 66,
  105, 66,
  106, 66,
  107, 66,
  108, 66,
  109, 66,
  110, 66,
  111, 66,
  112, 66,
  113, 66,
  114, 66,
  115, 66,
  116, 66,
  141, 66,
  142, 66,
  143, 66,
  144, 66,
  1, 67,
  2, 67,
  3, 67,
  4, 67,
  5, 67,
  6, 67,
  7, 67,
  8, 67,
  9, 67,
  10, 67,
  11, 67,
  12, 67,
  16, 67,
  17, 67,
  18, 67,
  19, 67,
  20, 67,
  21, 67,
  22, 67,
  23, 67,
  24, 67,
  25, 67,
  26, 67,
  27, 67,
  28, 67,
  29, 67,
  30, 67,
  31, 67,
  32, 67,
  33, 67,
  34, 67,
  35, 67,
  36, 67,
  37, 67,
  38, 67,
  39, 67,
  40, 67,
  41, 67,
  42, 67,
  43, 67,
  44, 67,
  45, 67,
  46, 67,
  47, 67,
  48, 67,
  49, 67,
  50, 67,
  51, 67,
  52, 67,
  53, 67,
  54, 67,
  55, 67,
  57, 67,
  58, 67,
  95, 67,
  96, 67,
  97, 67,
  98, 67,
  99, 67,
  100, 67,
  101, 67,
  102, 67,
  103, 67,
  104, 67,
  105, 67,
  106, 67,
  107, 67,
  108, 67,
  109, 67,
  110, 67,
  111, 67,
  112, 67,
  113, 67,
  114, 67,
  115, 67,
  116, 67,
  117, 67,
  118, 67,
  119, 67,
  141, 67,
  142, 67,
  143, 67,
  144, 67,
  1, 68,
  2, 68,
  3, 68,
  4, 68,
  5, 68,
  6, 68,
  7, 68,
  8, 68,
  9, 68,
  10, 68,
  11, 68,
  12, 68,
  13, 68,
  14, 68,
  15, 68,
  16, 68,
  17, 68,
  18, 68,
  19, 68,
  20, 68,
  21, 68,
  22, 68,
  23, 68,
  24, 68,
  25, 68,
  26, 68,
  27, 68,
  28, 68,
  29, 68,
  30, 68,
  31, 68,
  32, 68,
  33, 68,
  34, 68,
  35, 68,
  36, 68,
  37, 68,
  38, 68,
  39, 68,
  40, 68,
  41, 68,
  42, 68,
  43, 68,
  44, 68,
  45, 68,
  46, 68,
  47, 68,
  48, 68,
  49, 68,
  50, 68,
  51, 68,
  52, 68,
  53, 68,
  54, 68,
  55, 68,
  56, 68,
  57, 68,
  58, 68,
  95, 68,
  96, 68,
  97, 68,
  98, 68,
  99, 68,
  100, 68,
  101, 68,
  102, 68,
  103, 68,
  104, 68,
  105, 68,
  106, 68,
  107, 68,
  108, 68,
  109, 68,
  110, 68,
  111, 68,
  112, 68,
  113, 68,
  114, 68,
  115, 68,
  116, 68,
  117, 68,
  118, 68,
  119, 68,
  120, 68,
  144, 68,
  1, 69,
  2, 69,
  3, 69,
  4, 69,
  5, 69,
  6, 69,
  7, 69,
  8, 69,
  9, 69,
  10, 69,
  11, 69,
  12, 69,
  13, 69,
  14, 69,
  15, 69,
  16, 69,
  17, 69,
  18, 69,
  19, 69,
  20, 69,
  21, 69,
  22, 69,
  23, 69,
  24, 69,
  25, 69,
  26, 69,
  27, 69,
  28, 69,
  29, 69,
  30, 69,
  31, 69,
  32, 69,
  33, 69,
  34, 69,
  35, 69,
  36, 69,
  37, 69,
  38, 69,
  39, 69,
  40, 69,
  41, 69,
  42, 69,
  43, 69,
  44, 69,
  45, 69,
  46, 69,
  47, 69,
  48, 69,
  49, 69,
  50, 69,
  51, 69,
  52, 69,
  53, 69,
  54, 69,
  55, 69,
  56, 69,
  57, 69,
  58, 69,
  95, 69,
  96, 69,
  97, 69,
  98, 69,
  99, 69,
  100, 69,
  101, 69,
  102, 69,
  103, 69,
  104, 69,
  105, 69,
  106, 69,
  107, 69,
  108, 69,
  109, 69,
  110, 69,
  111, 69,
  112, 69,
  113, 69,
  114, 69,
  115, 69,
  116, 69,
  117, 69,
  118, 69,
  119, 69,
  121, 69,
  122, 69,
  123, 69,
  143, 69,
  144, 69,
  1, 70,
  2, 70,
  3, 70,
  4, 70,
  5, 70,
  6, 70,
  7, 70,
  8, 70,
  9, 70,
  10, 70,
  11, 70,
  12, 70,
  13, 70,
  14, 70,
  15, 70,
  16, 70,
  17, 70,
  18, 70,
  19, 70,
  20, 70,
  21, 70,
  22, 70,
  23, 70,
  24, 70,
  25, 70,
  26, 70,
  27, 70,
  28, 70,
  29, 70,
  30, 70,
  31, 70,
  32, 70,
  33, 70,
  34, 70,
  35, 70,
  36, 70,
  37, 70,
  38, 70,
  39, 70,
  40, 70,
  41, 70,
  42, 70,
  43, 70,
  44, 70,
  45, 70,
  46, 70,
  47, 70,
  48, 70,
  49, 70,
  50, 70,
  51, 70,
  52, 70,
  53, 70,
  54, 70,
  55, 70,
  56, 70,
  57, 70,
  58, 70,
  93, 70,
  94, 70,
  95, 70,
  96, 70,
  97, 70,
  98, 70,
  99, 70,
  100, 70,
  101, 70,
  102, 70,
  103, 70,
  104, 70,
  105, 70,
  106, 70,
  107, 70,
  108, 70,
  109, 70,
  110, 70,
  111, 70,
  112, 70,
  113, 70,
  114, 70,
  115, 70,
  116, 70,
  117, 70,
  118, 70,
  119, 70,
  120, 70,
  121, 70,
  122, 70,
  123, 70,
  143, 70,
  144, 70,
  1, 71,
  2, 71,
  3, 71,
  4, 71,
  5, 71,
  6, 71,
  7, 71,
  8, 71,
  9, 71,
  10, 71,
  11, 71,
  12, 71,
  13, 71,
  14, 71,
  15, 71,
  16, 71,
  17, 71,
  18, 71,
  19, 71,
  20, 71,
  21, 71,
  22, 71,
  23, 71,
  24, 71,
  25, 71,
  26, 71,
  27, 71,
  28, 71,
  29, 71,
  30, 71,
  31, 71,
  32, 71,
  33, 71,
  34, 71,
  35, 71,
  36, 71,
  37, 71,
  38, 71,
  39, 71,
  40, 71,
  41, 71,
  42, 71,
  43, 71,
  44, 71,
  45, 71,
  46, 71,
  47, 71,
  48, 71,
  49, 71,
  50, 71,
  51, 71,
  52, 71,
  53, 71,
  54, 71,
  55, 71,
  56, 71,
  57, 71,
  58, 71,
  63, 71,
  64, 71,
  93, 71,
  94, 71,
  95, 71,
  96, 71,
  97, 71,
  98, 71,
  99, 71,
  100, 71,
  101, 71,
  102, 71,
  103, 71,
  104, 71,
  105, 71,
  106, 71,
  107, 71,
  108, 71,
  109, 71,
  110, 71,
  111, 71,
  112, 71,
  113, 71,
  114, 71,
  115, 71,
  116, 71,
  117, 71,
  118, 71,
  119, 71,
  120, 71,
  121, 71,
  122, 71,
  141, 71,
  142, 71,
  143, 71,
  144, 71,
  1, 72,
  3, 72,
  4, 72,
  5, 72,
  6, 72,
  7, 72,
  8, 72,
  9, 72,
  10, 72,
  11, 72,
  12, 72,
  13, 72,
  14, 72,
  15, 72,
  16, 72,
  17, 72,
  18, 72,
  19, 72,
  20, 72,
  21, 72,
  22, 72,
  23, 72,
  24, 72,
  25, 72,
  26, 72,
  27, 72,
  28, 72,
  29, 72,
  30, 72,
  31, 72,
  32, 72,
  33, 72,
  34, 72,
  35, 72,
  36, 72,
  37, 72,
  38, 72,
  39, 72,
  40, 72,
  41, 72,
  42, 72,
  43, 72,
  44, 72,
  45, 72,
  46, 72,
  47, 72,
  48, 72,
  49, 72,
  50, 72,
  51, 72,
  52, 72,
  53, 72,
  54, 72,
  55, 72,
  56, 72,
  57, 72,
  58, 72,
  63, 72,
  64, 72,
  65, 72,
  77, 72,
  79, 72,
  92, 72,
  93, 72,
  94, 72,
  95, 72,
  96, 72,
  97, 72,
  98, 72,
  99, 72,
  100, 72,
  101, 72,
  102, 72,
  103, 72,
  104, 72,
  105, 72,
  106, 72,
  107, 72,
  108, 72,
  109, 72,
  110, 72,
  111, 72,
  112, 72,
  113, 72,
  114, 72,
  115, 72,
  116, 72,
  117, 72,
  118, 72,
  119, 72,
  120, 72,
  121, 72,
  122, 72,
  141, 72,
  142, 72,
  143, 72,
  144, 72,
  4, 73,
  5, 73,
  6, 73,
  7, 73,
  8, 73,
  9, 73,
  10, 73,
  11, 73,
  12, 73,
  13, 73,
  14, 73,
  15, 73,
  16, 73,
  17, 73,
  18, 73,
  19, 73,
  20, 73,
  21, 73,
  22, 73,
  23, 73,
  24, 73,
  25, 73,
  26, 73,
  27, 73,
  28, 73,
  29, 73,
  30, 73,
  31, 73,
  32, 73,
  33, 73,
  34, 73,
  35, 73,
  36, 73,
  37, 73,
  38, 73,
  39, 73,
  40, 73,
  41, 73,
  42, 73,
  43, 73,
  44, 73,
  45, 73,
  46, 73,
  47, 73,
  48, 73,
  49, 73,
  50, 73,
  51, 73,
  52, 73,
  53, 73,
  54, 73,
  55, 73,
  56, 73,
  63, 73,
  64, 73,
  65, 73,
  66, 73,
  79, 73,
  80, 73,
  81, 73,
  91, 73,
  92, 73,
  93, 73,
  94, 73,
  95, 73,
  96, 73,
  97, 73,
  98, 73,
  99, 73,
  100, 73,
  101, 73,
  102, 73,
  103, 73,
  104, 73,
  105, 73,
  106, 73,
  107, 73,
  108, 73,
  109, 73,
  110, 73,
  111, 73,
  112, 73,
  113, 73,
  114, 73,
  115, 73,
  116, 73,
  117, 73,
  118, 73,
  119, 73,
  120, 73,
  121, 73,
  122, 73,
  141, 73,
  142, 73,
  143, 73,
  144, 73,
  3, 74,
  4, 74,
  5, 74,
  6, 74,
  7, 74,
  9, 74,
  10, 74,
  11, 74,
  12, 74,
  13, 74,
  14, 74,
  15, 74,
  16, 74,
  17, 74,
  18, 74,
  19, 74,
  20, 74,
  21, 74,
  22, 74,
  23, 74,
  24, 74,
  25, 74,
  26, 74,
  27, 74,
  28, 74,
  29, 74,
  30, 74,
  31, 74,
  32, 74,
  33, 74,
  34, 74,
  35, 74,
  36, 74,
  37, 74,
  38, 74,
  39, 74,
  40, 74,
  41, 74,
  42, 74,
  43, 74,
  44, 74,
  45, 74,
  46, 74,
  47, 74,
  48, 74,
  49, 74,
  50, 74,
  51, 74,
  52, 74,
  53, 74,
  54, 74,
  55, 74,
  56, 74,
  57, 74,
  63, 74,
  64, 74,
  65, 74,
  66, 74,
  80, 74,
  81, 74,
  82, 74,
  83, 74,
  84, 74,
  89, 74,
  90, 74,
  91, 74,
  92, 74,
  93, 74,
  94, 74,
  95, 74,
  96, 74,
  97, 74,
  98, 74,
  99, 74,
  100, 74,
  101, 74,
  102, 74,
  103, 74,
  104, 74,
  105, 74,
  106, 74,
  107, 74,
  108, 74,
  109, 74,
  113, 74,
  114, 74,
  115, 74,
  116, 74,
  117, 74,
  118, 74,
  119, 74,
  120, 74,
  142, 74,
  143, 74,
  144, 74,
  3, 75,
  4, 75,
  5, 75,
  6, 75,
  7, 75,
  8, 75,
  9, 75,
  10, 75,
  11, 75,
  12, 75,
  13, 75,
  14, 75,
  15, 75,
  16, 75,
  17, 75,
  18, 75,
  19, 75,
  20, 75,
  21, 75,
  22, 75,
  23, 75,
  24, 75,
  25, 75,
  26, 75,
  27, 75,
  28, 75,
  29, 75,
  30, 75,
  31, 75,
  32, 75,
  33, 75,
  34, 75,
  35, 75,
  36, 75,
  37, 75,
  38, 75,
  39, 75,
  40, 75,
  41, 75,
  42, 75,
  43, 75,
  44, 75,
  45, 75,
  46, 75,
  47, 75,
  48, 75,
  49, 75,
  50, 75,
  51, 75,
  52, 75,
  53, 75,
  54, 75,
  55, 75,
  56, 75,
  57, 75,
  58, 75,
  59, 75,
  60, 75,
  61, 75,
  62, 75,
  64, 75,
  65, 75,
  66, 75,
  67, 75,
  68, 75,
  69, 75,
  78, 75,
  79, 75,
  80, 75,
  81, 75,
  82, 75,
  83, 75,
  84, 75,
  85, 75,
  86, 75,
  87, 75,
  88, 75,
  89, 75,
  90, 75,
  91, 75,
  92, 75,
  93, 75,
  94, 75,
  95, 75,
  96, 75,
  97, 75,
  98, 75,
  99, 75,
  100, 75,
  101, 75,
  102, 75,
  103, 75,
  104, 75,
  105, 75,
  106, 75,
  107, 75,
  113, 75,
  114, 75,
  115, 75,
  116, 75,
  117, 75,
  118, 75,
  119, 75,
  126, 75,
  127, 75,
  143, 75,
  144, 75,
  3, 76,
  4, 76,
  5, 76,
  6, 76,
  7, 76,
  8, 76,
  9, 76,
  10, 76,
  11, 76,
  12, 76,
  13, 76,
  14, 76,
  15, 76,
  16, 76,
  17, 76,
  18, 76,
  19, 76,
  20, 76,
  21, 76,
  22, 76,
  23, 76,
  24, 76,
  25, 76,
  26, 76,
  27, 76,
  28, 76,
  29, 76,
  30, 76,
  31, 76,
  32, 76,
  33, 76,
  34, 76,
  35, 76,
  36, 76,
  37, 76,
  38, 76,
  39, 76,
  40, 76,
  41, 76,
  42, 76,
  43, 76,
  44, 76,
  45, 76,
  46, 76,
  47, 76,
  48, 76,
  49, 76,
  50, 76,
  51, 76,
  52, 76,
  53, 76,
  54, 76,
  55, 76,
  56, 76,
  57, 76,
  58, 76,
  59, 76,
  60, 76,
  61, 76,
  62, 76,
  63, 76,
  64, 76,
  65, 76,
  66, 76,
  67, 76,
  68, 76,
  69, 76,
  70, 76,
  71, 76,
  72, 76,
  78, 76,
  79, 76,
  80, 76,
  81, 76,
  82, 76,
  83, 76,
  84, 76,
  85, 76,
  86, 76,
  87, 76,
  88, 76,
  89, 76,
  90, 76,
  91, 76,
  92, 76,
  93, 76,
  94, 76,
  95, 76,
  96, 76,
  97, 76,
  98, 76,
  99, 76,
  100, 76,
  101, 76,
  102, 76,
  103, 76,
  104, 76,
  105, 76,
  106, 76,
  107, 76,
  108, 76,
  113, 76,
  114, 76,
  115, 76,
  116, 76,
  117, 76,
  118, 76,
  125, 76,
  126, 76,
  127, 76,
  128, 76,
  141, 76,
  142, 76,
  144, 76,
  3, 77,
  4, 77,
  5, 77,
  6, 77,
  7, 77,
  8, 77,
  9, 77,
  10, 77,
  11, 77,
  12, 77,
  13, 77,
  14, 77,
  15, 77,
  16, 77,
  17, 77,
  18, 77,
  19, 77,
  20, 77,
  21, 77,
  22, 77,
  23, 77,
  24, 77,
  25, 77,
  26, 77,
  27, 77,
  28, 77,
  29, 77,
  30, 77,
  31, 77,
  32, 77,
  33, 77,
  34, 77,
  35, 77,
  36, 77,
  37, 77,
  38, 77,
  39, 77,
  40, 77,
  41, 77,
  42, 77,
  43, 77,
  44, 77,
  45, 77,
  46, 77,
  47, 77,
  48, 77,
  49, 77,
  50, 77,
  51, 77,
  52, 77,
  53, 77,
  54, 77,
  55, 77,
  56, 77,
  57, 77,
  58, 77,
  59, 77,
  60, 77,
  61, 77,
  62, 77,
  63, 77,
  64, 77,
  65, 77,
  66, 77,
  67, 77,
  68, 77,
  69, 77,
  70, 77,
  71, 77,
  72, 77,
  75, 77,
  76, 77,
  78, 77,
  79, 77,
  80, 77,
  81, 77,
  82, 77,
  83, 77,
  84, 77,
  85, 77,
  86, 77,
  87, 77,
  88, 77,
  89, 77,
  90, 77,
  91, 77,
  92, 77,
  93, 77,
  94, 77,
  95, 77,
  96, 77,
  97, 77,
  98, 77,
  99, 77,
  100, 77,
  101, 77,
  102, 77,
  103, 77,
  104, 77,
  105, 77,
  106, 77,
  107, 77,
  108, 77,
  109, 77,
  110, 77,
  111, 77,
  112, 77,
  113, 77,
  114, 77,
  115, 77,
  116, 77,
  117, 77,
  118, 77,
  119, 77,
  124, 77,
  125, 77,
  126, 77,
  127, 77,
  128, 77,
  136, 77,
  137, 77,
  138, 77,
  139, 77,
  141, 77,
  142, 77,
  5, 78,
  6, 78,
  7, 78,
  8, 78,
  9, 78,
  10, 78,
  11, 78,
  12, 78,
  13, 78,
  14, 78,
  15, 78,
  16, 78,
  17, 78,
  18, 78,
  19, 78,
  20, 78,
  21, 78,
  22, 78,
  23, 78,
  24, 78,
  25, 78,
  26, 78,
  27, 78,
  28, 78,
  29, 78,
  30, 78,
  31, 78,
  32, 78,
  33, 78,
  34, 78,
  35, 78,
  36, 78,
  37, 78,
  38, 78,
  39, 78,
  40, 78,
  41, 78,
  42, 78,
  43, 78,
  44, 78,
  45, 78,
  46, 78,
  47, 78,
  48, 78,
  49, 78,
  50, 78,
  51, 78,
  52, 78,
  53, 78,
  54, 78,
  55, 78,
  56, 78,
  57, 78,
  58, 78,
  59, 78,
  60, 78,
  61, 78,
  62, 78,
  63, 78,
  64, 78,
  65, 78,
  66, 78,
  67, 78,
  68, 78,
  69, 78,
  70, 78,
  71, 78,
  72, 78,
  73, 78,
  74, 78,
  75, 78,
  76, 78,
  77, 78,
  78, 78,
  79, 78,
  80, 78,
  81, 78,
  82, 78,
  83, 78,
  84, 78,
  85, 78,
  86, 78,
  87, 78,
  88, 78,
  89, 78,
  90, 78,
  91, 78,
  92, 78,
  93, 78,
  94, 78,
  95, 78,
  96, 78,
  97, 78,
  98, 78,
  99, 78,
  100, 78,
  101, 78,
  102, 78,
  103, 78,
  104, 78,
  105, 78,
  106, 78,
  107, 78,
  108, 78,
  109, 78,
  110, 78,
  111, 78,
  112, 78,
  113, 78,
  114, 78,
  115, 78,
  116, 78,
  117, 78,
  118, 78,
  119, 78,
  120, 78,
  123, 78,
  124, 78,
  125, 78,
  126, 78,
  127, 78,
  128, 78,
  129, 78,
  130, 78,
  131, 78,
  135, 78,
  136, 78,
  137, 78,
  138, 78,
  139, 78,
  6, 79,
  7, 79,
  8, 79,
  9, 79,
  10, 79,
  11, 79,
  12, 79,
  13, 79,
  14, 79,
  15, 79,
  16, 79,
  17, 79,
  18, 79,
  19, 79,
  20, 79,
  21, 79,
  22, 79,
  23, 79,
  24, 79,
  25, 79,
  26, 79,
  27, 79,
  28, 79,
  29, 79,
  30, 79,
  31, 79,
  32, 79,
  33, 79,
  34, 79,
  35, 79,
  36, 79,
  37, 79,
  38, 79,
  39, 79,
  40, 79,
  41, 79,
  42, 79,
  43, 79,
  44, 79,
  45, 79,
  46, 79,
  47, 79,
  48, 79,
  49, 79,
  50, 79,
  51, 79,
  52, 79,
  53, 79,
  54, 79,
  55, 79,
  56, 79,
  57, 79,
  58, 79,
  59, 79,
  60, 79,
  61, 79,
  62, 79,
  63, 79,
  64, 79,
  65, 79,
  66, 79,
  67, 79,
  68, 79,
  69, 79,
  70, 79,
  71, 79,
  72, 79,
  73, 79,
  74, 79,
  75, 79,
  76, 79,
  78, 79,
  79, 79,
  80, 79,
  81, 79,
  82, 79,
  83, 79,
  84, 79,
  85, 79,
  86, 79,
  87, 79,
  88, 79,
  89, 79,
  90, 79,
  91, 79,
  92, 79,
  93, 79,
  94, 79,
  95, 79,
  96, 79,
  97, 79,
  98, 79,
  99, 79,
  100, 79,
  101, 79,
  102, 79,
  103, 79,
  104, 79,
  105, 79,
  106, 79,
  107, 79,
  108, 79,
  109, 79,
  110, 79,
  111, 79,
  112, 79,
  114, 79,
  115, 79,
  116, 79,
  117, 79,
  118, 79,
  119, 79,
  120, 79,
  123, 79,
  124, 79,
  125, 79,
  126, 79,
  127, 79,
  128, 79,
  129, 79,
  130, 79,
  131, 79,
  132, 79,
  7, 80,
  8, 80,
  9, 80,
  10, 80,
  11, 80,
  12, 80,
  13, 80,
  14, 80,
  15, 80,
  16, 80,
  19, 80,
  20, 80,
  21, 80,
  22, 80,
  23, 80,
  24, 80,
  25, 80,
  26, 80,
  27, 80,
  28, 80,
  29, 80,
  30, 80,
  31, 80,
  32, 80,
  33, 80,
  34, 80,
  35, 80,
  36, 80,
  37, 80,
  38, 80,
  39, 80,
  40, 80,
  41, 80,
  42, 80,
  43, 80,
  44, 80,
  45, 80,
  46, 80,
  47, 80,
  48, 80,
  49, 80,
  50, 80,
  51, 80,
  52, 80,
  53, 80,
  54, 80,
  55, 80,
  56, 80,
  57, 80,
  58, 80,
  59, 80,
  60, 80,
  61, 80,
  62, 80,
  63, 80,
  64, 80,
  65, 80,
  66, 80,
  67, 80,
  68, 80,
  69, 80,
  70, 80,
  71, 80,
  72, 80,
  73, 80,
  78, 80,
  79, 80,
  80, 80,
  81, 80,
  82, 80,
  83, 80,
  84, 80,
  85, 80,
  86, 80,
  87, 80,
  88, 80,
  89, 80,
  90, 80,
  91, 80,
  92, 80,
  93, 80,
  94, 80,
  95, 80,
  96, 80,
  97, 80,
  98, 80,
  99, 80,
  100, 80,
  101, 80,
  102, 80,
  103, 80,
  104, 80,
  105, 80,
  106, 80,
  107, 80,
  108, 80,
  109, 80,
  110, 80,
  111, 80,
  112, 80,
  113, 80,
  114, 80,
  115, 80,
  116, 80,
  117, 80,
  118, 80,
  123, 80,
  124, 80,
  125, 80,
  126, 80,
  127, 80,
  128, 80,
  129, 80,
  130, 80,
  131, 80,
  132, 80,
  133, 80,
  134, 80,
  135, 80,
  9, 81,
  10, 81,
  11, 81,
  21, 81,
  22, 81,
  23, 81,
  27, 81,
  28, 81,
  29, 81,
  30, 81,
  31, 81,
  32, 81,
  33, 81,
  34, 81,
  35, 81,
  36, 81,
  37, 81,
  38, 81,
  39, 81,
  40, 81,
  41, 81,
  42, 81,
  43, 81,
  44, 81,
  45, 81,
  46, 81,
  47, 81,
  48, 81,
  49, 81,
  50, 81,
  51, 81,
  52, 81,
  53, 81,
  54, 81,
  55, 81,
  56, 81,
  57, 81,
  58, 81,
  59, 81,
  60, 81,
  61, 81,
  62, 81,
  63, 81,
  64, 81,
  72, 81,
  73, 81,
  81, 81,
  82, 81,
  83, 81,
  94, 81,
  95, 81,
  96, 81,
  97, 81,
  98, 81,
  99, 81,
  100, 81,
  101, 81,
  102, 81,
  103, 81,
  104, 81,
  105, 81,
  106, 81,
  107, 81,
  108, 81,
  109, 81,
  110, 81,
  111, 81,
  112, 81,
  113, 81,
  114, 81,
  115, 81,
  116, 81,
  117, 81,
  122, 81,
  123, 81,
  124, 81,
  125, 81,
  126, 81,
  127, 81,
  128, 81,
  129, 81,
  130, 81,
  131, 81,
  132, 81,
  133, 81,
  134, 81,
  135, 81,
  136, 81,
  21, 82,
  22, 82,
  23, 82,
  24, 82,
  28, 82,
  29, 82,
  30, 82,
  31, 82,
  32, 82,
  33, 82,
  34, 82,
  35, 82,
  36, 82,
  37, 82,
  38, 82,
  39, 82,
  40, 82,
  41, 82,
  42, 82,
  43, 82,
  44, 82,
  45, 82,
  46, 82,
  47, 82,
  48, 82,
  49, 82,
  50, 82,
  51, 82,
  52, 82,
  56, 82,
  57, 82,
  58, 82,
  59, 82,
  60, 82,
  61, 82,
  94, 82,
  95, 82,
  96, 82,
  97, 82,
  98, 82,
  99, 82,
  100, 82,
  101, 82,
  102, 82,
  103, 82,
  104, 82,
  105, 82,
  106, 82,
  107, 82,
  108, 82,
  109, 82,
  110, 82,
  111, 82,
  112, 82,
  113, 82,
  114, 82,
  122, 82,
  123, 82,
  124, 82,
  125, 82,
  126, 82,
  127, 82,
  128, 82,
  129, 82,
  130, 82,
  131, 82,
  132, 82,
  133, 82,
  134, 82,
  135, 82,
  136, 82,
  22, 83,
  23, 83,
  24, 83,
  25, 83,
  26, 83,
  27, 83,
  28, 83,
  35, 83,
  36, 83,
  37, 83,
  38, 83,
  39, 83,
  40, 83,
  41, 83,
  42, 83,
  43, 83,
  44, 83,
  45, 83,
  46, 83,
  47, 83,
  55, 83,
  56, 83,
  57, 83,
  58, 83,
  59, 83,
  60, 83,
  61, 83,
  95, 83,
  96, 83,
  97, 83,
  98, 83,
  99, 83,
  100, 83,
  101, 83,
  102, 83,
  103, 83,
  104, 83,
  105, 83,
  106, 83,
  107, 83,
  108, 83,
  109, 83,
  110, 83,
  111, 83,
  112, 83,
  113, 83,
  117, 83,
  118, 83,
  119, 83,
  120, 83,
  121, 83,
  122, 83,
  123, 83,
  124, 83,
  125, 83,
  126, 83,
  127, 83,
  128, 83,
  129, 83,
  130, 83,
  131, 83,
  132, 83,
  133, 83,
  134, 83,
  135, 83,
  136, 83,
  137, 83,
  5, 84,
  6, 84,
  7, 84,
  8, 84,
  9, 84,
  10, 84,
  26, 84,
  27, 84,
  39, 84,
  40, 84,
  41, 84,
  42, 84,
  43, 84,
  44, 84,
  45, 84,
  96, 84,
  97, 84,
  98, 84,
  99, 84,
  103, 84,
  104, 84,
  105, 84,
  106, 84,
  107, 84,
  108, 84,
  109, 84,
  110, 84,
  111, 84,
  112, 84,
  113, 84,
  114, 84,
  116, 84,
  117, 84,
  118, 84,
  119, 84,
  120, 84,
  121, 84,
  122, 84,
  123, 84,
  124, 84,
  125, 84,
  126, 84,
  127, 84,
  128, 84,
  129, 84,
  130, 84,
  131, 84,
  132, 84,
  133, 84,
  134, 84,
  135, 84,
  136, 84,
  137, 84,
  5, 85,
  6, 85,
  7, 85,
  8, 85,
  9, 85,
  10, 85,
  11, 85,
  12, 85,
  19, 85,
  20, 85,
  21, 85,
  22, 85,
  23, 85,
  24, 85,
  25, 85,
  26, 85,
  36, 85,
  37, 85,
  38, 85,
  39, 85,
  40, 85,
  41, 85,
  42, 85,
  43, 85,
  103, 85,
  104, 85,
  105, 85,
  106, 85,
  107, 85,
  108, 85,
  109, 85,
  110, 85,
  111, 85,
  112, 85,
  113, 85,
  114, 85,
  115, 85,
  116, 85,
  118, 85,
  119, 85,
  120, 85,
  121, 85,
  122, 85,
  123, 85,
  124, 85,
  125, 85,
  126, 85,
  127, 85,
  128, 85,
  129, 85,
  130, 85,
  131, 85,
  132, 85,
  133, 85,
  134, 85,
  135, 85,
  136, 85,
  137, 85,
  138, 85,
  20, 86,
  21, 86,
  22, 86,
  23, 86,
  25, 86,
  26, 86,
  37, 86,
  38, 86,
  39, 86,
  40, 86,
  107, 86,
  108, 86,
  109, 86,
  110, 86,
  111, 86,
  112, 86,
  113, 86,
  114, 86,
  115, 86,
  116, 86,
  117, 86,
  119, 86,
  120, 86,
  121, 86,
  122, 86,
  123, 86,
  124, 86,
  125, 86,
  126, 86,
  127, 86,
  128, 86,
  129, 86,
  130, 86,
  131, 86,
  132, 86,
  133, 86,
  134, 86,
  135, 86,
  136, 86,
  137, 86,
  138, 86,
  139, 86,
  111, 87,
  112, 87,
  113, 87,
  114, 87,
  115, 87,
  116, 87,
  117, 87,
  118, 87,
  127, 87,
  128, 87,
  129, 87,
  130, 87,
  131, 87,
  132, 87,
  133, 87,
  134, 87 ;

 xgrid_area = 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 275836070.864902, 275836070.864902, 275836070.864902, 
    275836070.864902, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 2206173067.44241, 2206173067.44241, 2206173067.44241, 
    2206173067.44241, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 4409597517.96414, 4409597517.96414, 4409597517.96414, 
    4409597517.96414, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 6607528159.0792, 6607528159.0792, 6607528159.0792, 
    6607528159.0792, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 6971823760.14062, 5429522593.37032, 
    5429522593.37032, 5429522593.37032, 5429522593.37032, 5429522593.37032, 
    5429522593.37032, 5429522593.37032, 5429522593.37032, 5429522593.37032, 
    5429522593.37032, 5429522593.37032, 5429522593.37032, 5429522593.37032, 
    5429522593.37032, 5429522593.37032, 10781708367.6144, 12119754811.1754, 
    12119754811.1754, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 12528264257.594, 
    12119754811.1754, 8105615480.49234, 5429522593.37032, 5429522593.37032, 
    5429522593.37032, 5429522593.37032, 5429522593.37032, 6767569036.93133, 
    12119754811.1754, 12324009534.3847, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 3600249646.33994, 6194612912.06638, 
    6194612912.06638, 6194612912.06638, 9290350035.85969, 13933955721.5497, 
    13933955721.5497, 14747414223.5798, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 14476261389.5697, 
    7742481473.96303, 2477845164.82645, 1238922582.41313, 6194612912.06638, 
    13933955721.5497, 15018567057.5899, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 14657491292.1255, 
    8758879986.09889, 1735660622.81716, 4142806465.20629, 6904677442.01039, 
    8660482282.83082, 15683701646.1126, 15683701646.1126, 15683701646.1126, 
    15683701646.1126, 15683701646.1126, 15683701646.1126, 15683701646.1126, 
    13927896805.2921, 6904677442.01039, 8660482282.83082, 17072230144.3662, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    15683701646.1126, 15683701646.1126, 15683701646.1126, 15683701646.1126, 
    16725098019.8028, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    2761870976.80424, 5523741953.60834, 12172091964.4717, 17072230144.3662, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    18231289940.5261, 17367281707.5436, 3923203884.01341, 6047417598.00796, 
    7559271997.50997, 7559271997.50997, 7559271997.50997, 7559271997.50997, 
    4535563198.50596, 16269687998.5194, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    6047417598.00796, 7559271997.50997, 15405679765.5369, 17367281707.5436, 
    17367281707.5436, 19527302289.9998, 19527302289.9998, 8158078602.51431, 
    8158078602.51431, 8158078602.51431, 8158078602.51431, 8158078602.51431, 
    8158078602.51431, 8158078602.51431, 8158078602.51431, 8158078602.51431, 
    8158078602.51431, 8158078602.51431, 12488096869.291, 18983124269.456, 
    21085355833.1183, 18983124269.456, 18983124269.456, 20559797942.2027, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 16818115136.0676, 
    8158078602.51431, 14653106002.6793, 21085355833.1183, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 18983124269.456, 18983124269.456, 8158078602.51431, 
    8158078602.51431, 3263231441.00578, 3263231441.00578, 10323087735.9026, 
    18983124269.456, 20559797942.2027, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 8158078602.51431, 8158078602.51431, 6960724224.44802, 
    5220543168.33602, 8700905280.56003, 15798241064.4647, 20529798253.7345, 
    23667600650.6441, 23667600650.6441, 23040040171.2622, 20529798253.7345, 
    20529798253.7345, 15798241064.4647, 8700905280.56002, 8700905280.56003, 
    6960724224.44802, 15798241064.4647, 20529798253.7345, 23667600650.6441, 
    22412479691.8803, 20529798253.7345, 21784919212.4984, 23667600650.6441, 
    23667600650.6441, 23667600650.6441, 23667600650.6441, 23667600650.6441, 
    23667600650.6441, 23667600650.6441, 23667600650.6441, 23040040171.2622, 
    20529798253.7345, 20529798253.7345, 20529798253.7345, 23040040171.2622, 
    20529798253.7345, 23667600650.6441, 23667600650.6441, 23667600650.6441, 
    21157358733.1165, 20529798253.7345, 20529798253.7345, 13432462469.8298, 
    8700905280.56003, 8700905280.56002, 8700905280.56003, 12317878952.2407, 
    21784919212.4984, 23667600650.6441, 23667600650.6441, 9187685618.91343, 
    9187685618.91343, 7350148495.13077, 9187685618.91343, 5512611371.3481, 
    3675074247.56543, 22006014214.3347, 22006014214.3347, 22006014214.3347, 
    11751351337.9977, 9187685618.91343, 9187685618.91343, 9187685618.91343, 
    9187685618.91343, 7350148495.13077, 7350148495.13077, 9187685618.91343, 
    9187685618.91343, 9187685618.91343, 1837537123.78277, 3675074247.56543, 
    19091954663.9816, 25694800694.027, 3688786479.69237, 737757295.938556, 
    5771086864.95806, 9618478108.26351, 17893766343.5355, 4682125033.40995, 
    1401293906.3744, 7006469531.87154, 7006469531.87154, 4203881719.12297, 
    20991196558.191, 37100304384.9128, 28760572874.4317, 6565970118.76537, 
    3425769697.09375, 38852825522.8721, 38852825522.8721, 15541130209.1488, 
    7696867319.82267, 15393734639.6454, 8029876190.72661, 16222776351.3347, 
    40556940878.3368, 40556940878.3368, 29883802977.645, 1877050145.19456, 
    8184944988.47009, 4438636545.67661, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 16795207361.5555, 4333075315.05564, 39382295100.9606, 
    13106159870.2092, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    17642323426.6722, 20958152656.1718, 2397902331.9947, 8757459419.42632, 
    33994039196.1925, 11678027494.0833, 31593492764.5643, 45357938424.7518, 
    45357938424.7518, 45357938424.7518, 33950527246.0276, 6790105449.2056, 
    11110111892.8723, 25529242158.8038, 10317851622.3745, 28108705064.3974, 
    46847841773.9957, 46847841773.9957, 46847841773.9957, 12897314527.9682, 
    2579462905.59371, 11056828790.3539, 11056828790.3539, 13783337023.25, 
    41387710034.4423, 2764207197.58847, 28967627127.6404, 48279378546.0673, 
    48279378546.0673, 48279378546.0673, 48279378546.0673, 20712704499.5673, 
    11056828790.3539, 39281080255.0127, 47576828230.5303, 47576828230.5303, 
    39281080255.0127, 5903288607.89877, 20178828463.5033, 2073936993.87941, 
    23887170526.7471, 49650765224.4097, 49650765224.4097, 49650765224.4097, 
    49650765224.4097, 49650765224.4097, 47576828230.5303, 7856216051.00256, 
    9423817467.4353, 9423817467.4353, 20739287584.3557, 40870988138.8763, 
    50960293231.9923, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    6282544978.29016, 24167422591.7669, 7050786157.25321, 47819020742.8472, 
    50960293231.9923, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    50960293231.9923, 22757148602.9789, 6282544978.29016, 33950907296.8275, 
    42438634121.0343, 42438634121.0343, 37283487434.846, 9997740414.05553, 
    31323798635.9911, 48299252284.4048, 42438634121.0343, 32128340748.6576, 
    6665160276.03706, 6665160276.03706, 52206331059.9851, 52206331059.9851, 
    52206331059.9851, 52206331059.9851, 52206331059.9851, 52206331059.9851, 
    27547692700.0311, 41765064847.9881, 52206331059.9851, 52206331059.9851, 
    52206331059.9851, 52206331059.9851, 52206331059.9851, 52206331059.9851, 
    41190566210.4263, 3332580138.01858, 3525046728.68103, 46234907769.0142, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 49624664200.8099, 
    7050093457.36213, 39082489237.612, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 47743333151.0067, 43980671051.4002, 43980671051.4002, 
    47743333151.0066, 53387326300.4164, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 51505995250.6131, 
    8796134210.27999, 42709861040.3331, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 35319827138.0055, 18344358794.4662, 54501807580.278, 
    54501807580.278, 54501807580.278, 54501807580.278, 54501807580.278, 
    29244720310.5218, 54501807580.278, 54501807580.278, 54501807580.278, 
    54501807580.278, 54501807580.278, 54501807580.278, 54501807580.278, 
    54501807580.278, 54501807580.278, 54501807580.278, 54501807580.278, 
    54501807580.278, 54501807580.278, 54501807580.278, 54501807580.278, 
    10900361516.0555, 36157448785.8117, 54501807580.278, 54501807580.278, 
    54501807580.278, 54501807580.278, 54501807580.278, 54501807580.278, 
    54501807580.278, 54501807580.278, 7443997278.41058, 52165407536.0034, 
    55548386394.6759, 55548386394.6759, 55548386394.6759, 55548386394.6759, 
    55548386394.6759, 53856896965.3396, 9418187849.59896, 18836375699.1979, 
    55548386394.6759, 55548386394.6759, 55548386394.6759, 55548386394.6759, 
    55548386394.6759, 55548386394.6759, 55548386394.6759, 55548386394.6759, 
    55548386394.6759, 55548386394.6759, 55548386394.6759, 55548386394.6759, 
    55548386394.6759, 55548386394.6759, 55548386394.6759, 11109677278.9352, 
    22219354557.8704, 55548386394.6759, 55548386394.6759, 55548386394.6759, 
    55548386394.6759, 55548386394.6759, 55548386394.6759, 55548386394.6759, 
    55548386394.6759, 41055730257.0682, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 29051101085.5377, 8872974659.09581, 28584813111.2532, 
    22610303534.692, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 52089271507.1822, 
    6868664437.7981, 22610303534.692, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 49657094398.932, 4436487329.5479, 
    21070385503.2943, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 33361742695.4771, 56481358529.3155, 10535192751.6471, 
    22973082888.8342, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 57432707222.0854, 57432707222.0854, 24875780274.3741, 
    1902697385.53996, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 57432707222.0854, 53627312451.0056, 25971649516.6072, 
    5194329903.32147, 36030882286.3438, 58268101605.9897, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 58268101605.9897, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 33890839640.8439, 58268101605.9897, 
    14132981902.7119, 10244280062.4339, 170987443.908059, 41825417589.7709, 
    54549059233.7188, 58268101605.9897, 58268101605.9897, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 58268101605.9897, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 58268101605.9897, 58268101605.9897, 
    43065098380.5279, 170987443.90806, 10412611554.54, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 58268101605.9897, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 58268101605.9897, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 37269235101.1998, 8016498943.22077, 
    55241219896.0749, 59030901191.0676, 59030901191.0676, 59030901191.0676, 
    59030901191.0676, 59030901191.0676, 59030901191.0676, 59030901191.0676, 
    59030901191.0676, 22205655839.4525, 23612360476.4271, 59030901191.0676, 
    35418540714.6406, 7579362589.98562, 36825245351.6152, 59030901191.0676, 
    59030901191.0676, 59030901191.0676, 59030901191.0676, 59030901191.0676, 
    59030901191.0676, 59030901191.0676, 59030901191.0676, 59030901191.0676, 
    44841744294.836, 3789681294.99283, 59030901191.0676, 59030901191.0676, 
    59030901191.0676, 59030901191.0676, 59030901191.0676, 59030901191.0676, 
    59030901191.0676, 59030901191.0676, 59030901191.0676, 59030901191.0676, 
    59030901191.0676, 59030901191.0676, 11944031124.8045, 59720155624.0228, 
    59720155624.0228, 59720155624.0228, 59720155624.0228, 59720155624.0228, 
    59720155624.0228, 59720155624.0228, 59720155624.0228, 59720155624.0228, 
    53257735702.2698, 27408056015.2578, 12924839843.506, 57992035648.2724, 
    56239057009.8566, 6462419921.75296, 43275322014.8681, 59720155624.0228, 
    59720155624.0228, 59720155624.0228, 59720155624.0228, 58856095636.1476, 
    36929650823.9413, 47028813242.1693, 59720155624.0228, 23888062249.6091, 
    4721870614.66987, 13956973045.0226, 7209731178.80197, 36851797244.5976, 
    59720155624.0228, 59720155624.0228, 59720155624.0228, 59720155624.0228, 
    59720155624.0228, 59720155624.0228, 59720155624.0228, 59720155624.0228, 
    59720155624.0228, 59720155624.0228, 59720155624.0228, 59720155624.0228, 
    20406963635.4429, 12067001235.9321, 60335006179.6604, 60335006179.6604, 
    60335006179.6604, 60335006179.6604, 60335006179.6604, 60335006179.6604, 
    60335006179.6604, 60335006179.6604, 60335006179.6604, 60335006179.6604, 
    60335006179.6604, 15377123559.0006, 56340654138.3353, 7304474364.39368, 
    60335006179.6604, 60335006179.6604, 60335006179.6604, 60335006179.6604, 
    31438476836.2578, 12067001235.9321, 60335006179.6604, 7304474364.39367, 
    16829528107.4705, 53030531815.2667, 60335006179.6604, 60335006179.6604, 
    60335006179.6604, 60335006179.6604, 60335006179.6604, 60335006179.6604, 
    60335006179.6604, 60335006179.6604, 60335006179.6604, 60335006179.6604, 
    60335006179.6604, 60335006179.6604, 60335006179.6604, 24134002471.8642, 
    337729666.551555, 49037479131.1532, 60874686830.752, 60874686830.752, 
    60874686830.752, 60874686830.752, 60874686830.752, 60874686830.752, 
    60874686830.752, 60874686830.752, 60874686830.752, 60874686830.752, 
    26736254145.4621, 1688648332.7578, 1688648332.75779, 60874686830.752, 
    60874686830.752, 39517622579.2026, 12174937366.1504, 30404523959.3166, 
    39517622579.2026, 60874686830.752, 60874686830.752, 60874686830.752, 
    60874686830.752, 60874686830.752, 60874686830.752, 60874686830.752, 
    60874686830.752, 60874686830.752, 60874686830.752, 60874686830.752, 
    60874686830.752, 60874686830.752, 60874686830.752, 31145622204.5386, 
    49070820161.9277, 61338525202.4097, 61338525202.4097, 61338525202.4097, 
    61338525202.4097, 61338525202.4097, 61338525202.4097, 61338525202.4097, 
    61338525202.4097, 61338525202.4097, 61338525202.4097, 6749889103.53542, 
    11852521903.3458, 3669054035.92654, 2935243228.74122, 12267705040.4819, 
    12267705040.4819, 6749889103.53542, 7442160299.58697, 56512980461.5147, 
    61338525202.4097, 61338525202.4097, 61338525202.4097, 61338525202.4097, 
    61338525202.4097, 61338525202.4097, 61338525202.4097, 61338525202.4097, 
    61338525202.4097, 61338525202.4097, 61338525202.4097, 61338525202.4097, 
    61338525202.4097, 61338525202.4097, 60604714395.2243, 18283783336.832, 
    49380754727.8242, 61725943409.7802, 61725943409.7802, 61725943409.7802, 
    61725943409.7802, 61725943409.7802, 61725943409.7802, 61725943409.7802, 
    61725943409.7802, 61725943409.7802, 46516749877.3188, 10695397026.0355, 
    25904590558.497, 14260529368.0474, 17560112679.8884, 8078928848.43772, 
    27554382214.4175, 12345188681.956, 18791498289.6714, 35966709811.7536, 
    1367910152.61661, 27554382214.4175, 61725943409.7802, 61725943409.7802, 
    61725943409.7802, 61725943409.7802, 61725943409.7802, 61725943409.7802, 
    61725943409.7802, 61725943409.7802, 61725943409.7802, 61725943409.7802, 
    61725943409.7802, 61725943409.7802, 61725943409.7802, 61725943409.7802, 
    61725943409.7802, 61725943409.7802, 52244759578.3295, 4201300721.63807, 
    53830467744.055, 62036458778.0211, 62036458778.0211, 62036458778.0211, 
    62036458778.0211, 62036458778.0211, 62036458778.0211, 62036458778.0211, 
    62036458778.0211, 62036458778.0211, 37221875266.8127, 27596334224.1196, 
    50072482278.1467, 38869300281.9855, 23321580169.1913, 1296392932.70716, 
    2160654887.84526, 1728523910.27621, 7862241387.06824, 933813445.835339, 
    47900643112.1407, 61172196822.883, 60307934867.7449, 52931430043.5683, 
    5100338422.12479, 933813445.835341, 7468787997.44079, 933813445.835339, 
    61172196822.883, 62036458778.0211, 62036458778.0211, 62036458778.0211, 
    62036458778.0211, 62036458778.0211, 62036458778.0211, 62036458778.0211, 
    62036458778.0211, 62036458778.0211, 62036458778.0211, 62036458778.0211, 
    62036458778.0211, 62036458778.0211, 62036458778.0211, 62036458778.0211, 
    62036458778.0211, 62036458778.0211, 17500002986.1659, 62269684443.65, 
    62269684443.65, 62269684443.65, 62269684443.65, 62269684443.65, 
    62269684443.65, 62269684443.65, 62269684443.65, 62269684443.65, 
    62269684443.65, 42407876763.6259, 2523033048.71796, 32832131650.5203, 
    24907873777.46, 18623944816.7864, 15934709087.3798, 5842576892.50801, 
    11329995058.1096, 29212884462.54, 55658324447.428, 62269684443.65, 
    57223618346.2141, 19506648953.1177, 6283928960.67369, 13222719992.444, 
    24907873777.46, 62269684443.65, 62269684443.65, 62269684443.65, 
    62269684443.65, 62269684443.65, 62269684443.65, 62269684443.65, 
    62269684443.65, 62269684443.65, 62269684443.65, 62269684443.65, 
    62269684443.65, 62269684443.65, 62269684443.65, 62269684443.65, 
    62269684443.65, 56427107551.142, 33056799981.1101, 1493851821.06265, 
    55136673902.0721, 62425329836.5296, 62425329836.5296, 62425329836.5296, 
    62425329836.5296, 62425329836.5296, 62425329836.5296, 62425329836.5296, 
    62425329836.5296, 62425329836.5296, 62425329836.5296, 62425329836.5296, 
    1493851821.06265, 19083362659.4216, 62425329836.5296, 41157756113.7036, 
    32816619993.5905, 44203690000.386, 23689895843.335, 24970131934.6118, 
    50580381914.8621, 640118045.638437, 6008419843.18056, 22166358616.0774, 
    14849157843.2578, 56006913956.9613, 60931478015.4669, 60931478015.4669, 
    40387998452.221, 4924564058.50559, 7878532783.39257, 62425329836.5296, 
    62425329836.5296, 62425329836.5296, 62425329836.5296, 62425329836.5296, 
    62425329836.5296, 62425329836.5296, 62425329836.5296, 62425329836.5296, 
    62425329836.5296, 62425329836.5296, 62425329836.5296, 62425329836.5296, 
    62425329836.5296, 56138477848.3464, 45929588106.2403, 8568892025.73431, 
    25001280416.7528, 62503201041.8819, 62503201041.8819, 62503201041.8819, 
    62503201041.8819, 62503201041.8819, 62503201041.8819, 62503201041.8819, 
    62503201041.8819, 62503201041.8819, 62503201041.8819, 62503201041.8819, 
    62503201041.8819, 44100044258.721, 2067046925.10773, 54533637541.9897, 
    49901028163.7009, 3351290509.02905, 17031716916.8605, 62503201041.8819, 
    62503201041.8819, 46651270324.4765, 7969563499.89221, 46040702609.5618, 
    8974892555.16878, 6468375389.55624, 6468375389.55624, 19146832411.8799, 
    27116395911.7721, 5026935763.54358, 5026935763.54358, 16682802628.5034, 
    62503201041.8819, 62503201041.8819, 62503201041.8819, 62503201041.8819, 
    62503201041.8819, 62503201041.8819, 62503201041.8819, 62503201041.8819, 
    62503201041.8819, 62503201041.8819, 62503201041.8819, 58369107191.6664, 
    45891390509.2924, 24280528314.0361, 17031726805.4509, 62503201041.8819, 
    62503201041.8819, 62503201041.8819, 62503201041.8819, 62503201041.8819, 
    62503201041.8819, 62503201041.8819, 62503201041.8819, 62503201041.8819, 
    62503201041.8819, 62503201041.8819, 62503201041.8819, 62503201041.8819, 
    32534713568.3122, 4356619563.21705, 41906588976.2094, 62503201041.8819, 
    28788681498.695, 25001280416.7527, 62503201041.8819, 62503201041.8819, 
    58343957202.3735, 8341396368.86799, 18878758674.3457, 14989815032.7146, 
    10824999897.2764, 27507792635.0124, 42469127681.946, 62503201041.8819, 
    62503201041.8819, 62503201041.8819, 62503201041.8819, 62503201041.8819, 
    62503201041.8819, 62503201041.8819, 62503201041.8819, 62503201041.8819, 
    62503201041.8819, 55017816678.1856, 1280226223.21903, 62425329836.5296, 
    62425329836.5296, 62425329836.5296, 62425329836.5296, 62425329836.5296, 
    62425329836.5296, 62425329836.5296, 62425329836.5296, 62425329836.5296, 
    62425329836.5296, 62425329836.5296, 62425329836.5296, 62425329836.5296, 
    62425329836.5296, 31405029401.6075, 640113111.609516, 10466138903.665, 
    50557304265.4727, 55136683775.5517, 30166551840.9399, 1493861705.59169, 
    6286876698.04337, 51959190932.8646, 62425329836.5296, 12485065967.3059, 
    1493861705.59169, 8840742936.81699, 58781006806.0406, 62425329836.5296, 
    62425329836.5296, 62425329836.5296, 62425329836.5296, 62425329836.5296, 
    62425329836.5296, 62425329836.5296, 62425329836.5296, 62425329836.5296, 
    36174971678.6987, 6283919115.70318, 43015406866.2029, 54700570505.134, 
    62269684443.65, 62269684443.65, 62269684443.65, 62269684443.65, 
    62269684443.65, 62269684443.65, 62269684443.65, 62269684443.65, 
    62269684443.65, 62269684443.65, 62269684443.65, 62269684443.65, 
    62269684443.65, 62269684443.65, 62269684443.65, 25676647027.2589, 
    31405327504.0481, 5842581819.46556, 50584520804.7189, 12453936888.73, 
    11685163638.9311, 55985765327.9469, 26031815591.4762, 6283919115.70318, 
    49815747554.92, 62269684443.65, 62269684443.65, 62269684443.65, 
    62269684443.65, 62269684443.65, 62269684443.65, 62269684443.65, 
    55985765327.9469, 43090491142.9792, 5842581819.46556, 36376319186.2825, 
    36376319186.2825, 33056775346.3223, 26117984323.4965, 60635723857.3006, 
    59701900576.8203, 62036458778.0211, 62036458778.0211, 62036458778.0211, 
    62036458778.0211, 62036458778.0211, 62036458778.0211, 62036458778.0211, 
    62036458778.0211, 62036458778.0211, 62036458778.0211, 62036458778.0211, 
    62036458778.0211, 62036458778.0211, 62036458778.0211, 62036458778.0211, 
    62036458778.0211, 62036458778.0211, 45948368799.4571, 432126080.207836, 
    432126080.207845, 46897268301.0406, 9590745693.06011, 32819854257.1695, 
    466911640.240174, 13036042979.4127, 4633431713.27613, 3931120686.11437, 
    36538374449.4869, 32676824883.4372, 432126080.207836, 10022871773.2679, 
    9934490443.36729, 57835153144.9528, 62036458778.0211, 62036458778.0211, 
    62036458778.0211, 62036458778.0211, 62036458778.0211, 62036458778.0211, 
    36554248249.9977, 5135128913.54863, 432126080.207836, 40724858556.0078, 
    62036458778.0211, 62036458778.0211, 62036458778.0211, 62036458778.0211, 
    61725943409.7802, 61725943409.7802, 61725943409.7802, 61725943409.7802, 
    61725943409.7802, 61725943409.7802, 61725943409.7802, 61725943409.7802, 
    61725943409.7802, 61725943409.7802, 61725943409.7802, 61725943409.7802, 
    61725943409.7802, 61725943409.7802, 61725943409.7802, 61725943409.7802, 
    61725943409.7802, 61725943409.7802, 61725943409.7802, 61725943409.7802, 
    17560102901.5418, 21826362752.9337, 31307536823.9113, 15209203292.9345, 
    39899580656.8465, 1367900411.44054, 19611953518.7026, 683950205.720274, 
    7604601646.46723, 17085775717.4448, 33188552237.7228, 15209203292.9345, 
    1367900411.44054, 34645878618.9867, 38023008232.3362, 42096817476.5911, 
    34017888646.0269, 61725943409.7802, 61725943409.7802, 61725943409.7802, 
    60358042998.3397, 60358042998.3397, 44165840508.2383, 23194263164.3742, 
    61725943409.7802, 61725943409.7802, 61725943409.7802, 61725943409.7802, 
    61725943409.7802, 61338525202.4097, 61338525202.4097, 61338525202.4097, 
    61338525202.4097, 61338525202.4097, 61338525202.4097, 61338525202.4097, 
    61338525202.4097, 61338525202.4097, 61338525202.4097, 61338525202.4097, 
    61338525202.4097, 61338525202.4097, 61338525202.4097, 61338525202.4097, 
    61338525202.4097, 61338525202.4097, 33901934162.1265, 20941962796.8886, 
    37210825744.0008, 23067798141.4077, 38270727061.0019, 61338525202.4097, 
    42320921337.8835, 733805969.778028, 43054727307.6616, 61338525202.4097, 
    30053216297.4016, 14884330297.6003, 8158949658.68173, 57229769820.6095, 
    26003022020.52, 31285308905.0081, 33168128192.3484, 41302559665.9045, 
    41327077851.0302, 10124848236.0663, 10124848236.0663, 10124848236.0663, 
    2935223879.1122, 61338525202.4097, 61338525202.4097, 61338525202.4097, 
    61338525202.4097, 61338525202.4097, 61338525202.4097, 60874686830.752, 
    60874686830.752, 60874686830.752, 60874686830.752, 60874686830.752, 
    60874686830.752, 60874686830.752, 60874686830.752, 60874686830.752, 
    60874686830.752, 60874686830.752, 60874686830.752, 60874686830.752, 
    60874686830.752, 60874686830.752, 60874686830.752, 59861512221.1961, 
    46945447717.3429, 18701959395.7373, 1013174609.55589, 675449739.703929, 
    60874686830.752, 60874686830.752, 48699749464.6016, 47283172587.1948, 
    60874686830.752, 60874686830.752, 36524812098.4512, 14110900764.2659, 
    34723515875.9949, 1350899479.40785, 22955293157.3566, 53290808096.0729, 
    41903992342.823, 48699749464.6016, 60874686830.752, 60874686830.752, 
    60874686830.752, 60874686830.752, 60874686830.752, 60874686830.752, 
    60335006179.6604, 60335006179.6604, 60335006179.6604, 60335006179.6604, 
    60335006179.6604, 60335006179.6604, 60335006179.6604, 60335006179.6604, 
    60335006179.6604, 60335006179.6604, 60335006179.6604, 60335006179.6604, 
    60335006179.6604, 60335006179.6604, 60335006179.6604, 53030541343.9366, 
    7988713644.84704, 48268004943.7283, 60335006179.6604, 52346292534.8134, 
    23449753662.7409, 31438467307.5879, 60335006179.6604, 60335006179.6604, 
    7304464835.7238, 48268004943.7283, 60335006179.6604, 60335006179.6604, 
    60335006179.6604, 28896538872.0725, 48268004943.7283, 3652232417.86191, 
    18261162089.3095, 22681574084.9562, 56340649357.2369, 56682773761.7985, 
    42073844090.3509, 33659075272.2807, 40963540108.0045, 60335006179.6604, 
    60335006179.6604, 60335006179.6604, 60335006179.6604, 60335006179.6604, 
    60335006179.6604, 59720155624.0228, 59720155624.0228, 59720155624.0228, 
    59720155624.0228, 59720155624.0228, 59720155624.0228, 59720155624.0228, 
    59720155624.0228, 59720155624.0228, 59720155624.0228, 59720155624.0228, 
    59720155624.0228, 59720155624.0228, 59720155624.0228, 59720155624.0228, 
    32351004172.5704, 9943504396.63999, 54238539694.015, 59720155624.0228, 
    59720155624.0228, 58856090889.8297, 36929627169.7985, 6962178403.6865, 
    47776124499.2182, 59720155624.0228, 59720155624.0228, 52510410225.6289, 
    9943504396.63999, 22159932781.2229, 41547178365.6133, 54238539694.015, 
    59720155624.0228, 59720155624.0228, 45159100031.568, 4345153936.0363, 
    40813946095.5317, 5221633802.76486, 18146464192.3584, 47028794295.6211, 
    59720155624.0228, 51017432619.4146, 57979611023.1012, 47776124499.2182, 
    1740544600.92158, 8702723004.60814, 3481089201.84322, 23888062249.6091, 
    59720155624.0228, 59720155624.0228, 59720155624.0228, 59720155624.0228, 
    59720155624.0228, 59720155624.0228, 59030901191.0676, 59030901191.0676, 
    59030901191.0676, 59030901191.0676, 59030901191.0676, 59030901191.0676, 
    59030901191.0676, 59030901191.0676, 59030901191.0676, 59030901191.0676, 
    59030901191.0676, 59030901191.0676, 59030901191.0676, 59030901191.0676, 
    50311054613.2094, 3086333660.3553, 42997893984.7378, 59030901191.0676, 
    59030901191.0676, 59030901191.0676, 59030901191.0676, 59030901191.0676, 
    55944567530.7124, 8719846577.8583, 47224720952.8541, 59030901191.0676, 
    59030901191.0676, 59030901191.0676, 52858233870.3571, 7579353270.09724, 
    31191713746.5243, 59030901191.0676, 59030901191.0676, 59030901191.0676, 
    59030901191.0676, 23612360476.4271, 16033007206.3299, 17439693155.7166, 
    7579353270.09724, 42997893984.7378, 59030901191.0676, 59030901191.0676, 
    34011854765.2539, 22205674527.0404, 47224720952.8541, 15158706540.1944, 
    8016503603.16496, 40082518015.8246, 9860339885.61937, 6172667320.71055, 
    23612360476.4271, 59030901191.0676, 59030901191.0676, 59030901191.0676, 
    59030901191.0676, 59030901191.0676, 59030901191.0676, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 58268101605.9897, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 58268101605.9897, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 58268101605.9897, 58268101605.9897, 
    58268101605.9897, 46614481284.7918, 20827869792.1276, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 58268101605.9897, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 43065079897.5882, 10583589784.2626, 
    52069674480.319, 57028416180.8556, 58268101605.9897, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 49426905326.6548, 16046362964.2052, 
    10755891471.6862, 57028416180.8556, 58268101605.9897, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 49426905326.6548, 26458974460.6566, 
    39182625318.7899, 5633751467.75369, 170978287.81118, 2479370850.26831, 
    10583589784.2626, 58268101605.9897, 58268101605.9897, 52976306713.8584, 
    6361825429.06661, 25447301716.2665, 256467431.716774, 427445719.527961, 
    31324647032.8723, 25531467460.5597, 43964132146.7123, 58268101605.9897, 
    58268101605.9897, 58268101605.9897, 58268101605.9897, 58268101605.9897, 
    58268101605.9897, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 57432707222.0854, 57432707222.0854, 52238372771.546, 
    41849703870.4672, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 56481363043.9078, 54578674687.5526, 56481363043.9078, 
    31312535068.3971, 951344178.177638, 36508841054.7671, 57432707222.0854, 
    57432707222.0854, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 26120172153.6883, 951344178.177638, 33654808520.2343, 
    12584413987.7554, 951344178.177638, 36508841054.7671, 57432707222.0854, 
    57432707222.0854, 45946165777.6683, 15583003351.6183, 25971672252.6971, 
    10388668901.0788, 21070394532.4789, 57432707222.0854, 57432707222.0854, 
    57432707222.0854, 57432707222.0854, 57432707222.0854, 57432707222.0854, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    45220607069.3841, 8872983619.45909, 32932515251.4026, 7246140486.25736, 
    34343299788.0824, 34343299788.0824, 38779791597.8119, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 25042471682.579, 
    8872983619.45908, 1449228097.25145, 21161075437.4406, 14203607961.849, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 46669835166.6356, 
    1449228097.25146, 5796912389.00589, 53627302642.2272, 56525758836.7301, 
    56525758836.7301, 56525758836.7301, 56525758836.7301, 56525758836.7301, 
    55548386394.6756, 55548386394.6756, 55548386394.6756, 55548386394.6756, 
    55548386394.6756, 55548386394.6756, 55548386394.6756, 55548386394.6756, 
    55548386394.6756, 55548386394.6756, 55548386394.6756, 55548386394.6756, 
    55548386394.6756, 55548386394.6756, 55548386394.6756, 55548386394.6756, 
    55548386394.6756, 55548386394.6756, 55548386394.6756, 55548386394.6756, 
    51562972748.698, 35621318164.7876, 47577559102.7204, 55548386394.6756, 
    55548386394.6756, 55548386394.6756, 55548386394.6756, 55548386394.6756, 
    55548386394.6756, 55548386394.6756, 55548386394.6756, 55548386394.6756, 
    55548386394.6756, 55548386394.6756, 55548386394.6756, 55548386394.6756, 
    55548386394.6756, 55548386394.6756, 55548386394.6756, 55548386394.6756, 
    55548386394.6756, 55548386394.6756, 55548386394.6756, 55548386394.6756, 
    55548386394.6756, 55548386394.6756, 55548386394.6756, 47577559102.7204, 
    17631497391.3018, 25358204544.8501, 17875617529.7086, 47577559102.7204, 
    55548386394.6756, 55548386394.6756, 55548386394.6756, 55548386394.6756, 
    11109677278.9351, 7124263632.95747, 48180002623.3112, 17389019508.1969, 
    50473931206.5955, 55548386394.6756, 55548386394.6756, 55548386394.6756, 
    55548386394.6756, 54501807580.2781, 54501807580.2781, 54501807580.2781, 
    54501807580.2781, 54501807580.2781, 54501807580.2781, 54501807580.2781, 
    54501807580.2781, 54501807580.2781, 54501807580.2781, 54501807580.2781, 
    54501807580.2781, 54501807580.2781, 54501807580.2781, 54501807580.2781, 
    54501807580.2781, 54501807580.2781, 54501807580.2781, 54501807580.2781, 
    54501807580.2781, 54501807580.2781, 54501807580.2781, 54501807580.2781, 
    54501807580.2781, 54501807580.2781, 54501807580.2781, 54501807580.2781, 
    54501807580.2781, 54501807580.2781, 54501807580.2781, 54501807580.2781, 
    54501807580.2781, 54501807580.2781, 54501807580.2781, 54501807580.2781, 
    54501807580.2781, 54501807580.2781, 54501807580.2781, 54501807580.2781, 
    54501807580.2781, 54501807580.2781, 54501807580.2781, 54501807580.2781, 
    54501807580.2781, 54501807580.2781, 54501807580.2781, 54501807580.2781, 
    54501807580.2781, 43601446064.2225, 3603214278.52554, 47057801650.6704, 
    54501807580.2781, 54501807580.2781, 54501807580.2781, 54501807580.2781, 
    54501807580.2781, 54501807580.2781, 39613795721.0628, 35891792756.259, 
    35891792756.259, 19761538520.2919, 9008035696.31381, 18106790073.1067, 
    32701084548.1668, 7444005929.60763, 54501807580.2781, 54501807580.2781, 
    54501807580.2781, 54501807580.2781, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 53387326300.4164, 
    28167429712.969, 17625254839.9733, 53387326300.4164, 45862018878.0533, 
    17625254839.9732, 17625254839.9733, 38709604585.9647, 28167429712.969, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 53387326300.4164, 38947207329.1516, 18067482295.3587, 
    35659759104.3438, 53387326300.4164, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 53387326300.4164, 
    53387326300.4164, 53387326300.4164, 35795049491.4313, 49624672589.2348, 
    53387326300.4164, 53387326300.4164, 53387326300.4164, 52206331059.9855, 
    52206331059.9855, 52206331059.9855, 52206331059.9855, 30880285281.5511, 
    16662921429.2614, 16662921429.2614, 3332584285.85239, 48299260484.7883, 
    52206331059.9855, 52206331059.9855, 52206331059.9855, 52206331059.9855, 
    52206331059.9855, 52206331059.9855, 52206331059.9855, 52206331059.9855, 
    52206331059.9855, 52206331059.9855, 52206331059.9855, 52206331059.9855, 
    52206331059.9855, 52206331059.9855, 52206331059.9855, 52206331059.9855, 
    52206331059.9855, 52206331059.9855, 52206331059.9855, 52206331059.9855, 
    52206331059.9855, 52206331059.9855, 52206331059.9855, 52206331059.9855, 
    52206331059.9855, 52206331059.9855, 52206331059.9855, 52206331059.9855, 
    52206331059.9855, 52206331059.9855, 52206331059.9855, 52206331059.9855, 
    52206331059.9855, 16975461848.797, 3907070575.19739, 34656382921.8436, 
    25233116353.6318, 7814141150.39464, 14922823076.5395, 48873746774.1333, 
    52206331059.9855, 52206331059.9855, 52206331059.9855, 52206331059.9855, 
    52206331059.9855, 52206331059.9855, 52206331059.9855, 52206331059.9855, 
    52206331059.9855, 52206331059.9855, 52206331059.9855, 52206331059.9855, 
    52206331059.9855, 52206331059.9855, 20077969715.0856, 1953535287.59877, 
    15152899496.1031, 46345725197.1896, 52206331059.9855, 52206331059.9855, 
    42888865162.2007, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    20384117292.7969, 4035714034.8957, 10089285087.2394, 6053571052.34361, 
    30576175939.1953, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    50960293231.9923, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    50960293231.9923, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    50960293231.9923, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    50960293231.9923, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    50960293231.9923, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    50960293231.9923, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    50960293231.9923, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    50960293231.9923, 50960293231.9923, 4035714034.8957, 27434899398.7497, 
    21152346317.8583, 9423829621.3369, 35838083056.2479, 43783302656.6508, 
    35253910529.7639, 4035714034.8957, 18137278246.8013, 50960293231.9923, 
    50960293231.9923, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    50960293231.9923, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    50960293231.9923, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    50960293231.9923, 50960293231.9923, 50960293231.9923, 50960293231.9923, 
    24293622858.304, 20384117292.7969, 15706382702.2283, 15706382702.2283, 
    2951648253.78075, 14758241268.9036, 14758241268.9036, 14758241268.9036, 
    5903296507.56147, 19618286778.0243, 4147866193.1903, 11126370984.2915, 
    11126370984.2915, 11126370984.2915, 40795820463.0675, 49650765224.4097, 
    43747468716.8482, 43747468716.8482, 49650765224.4097, 49650765224.4097, 
    49650765224.4097, 49650765224.4097, 49650765224.4097, 49650765224.4097, 
    49650765224.4097, 49650765224.4097, 49650765224.4097, 49650765224.4097, 
    49650765224.4097, 49650765224.4097, 49650765224.4097, 49650765224.4097, 
    49650765224.4097, 49650765224.4097, 49650765224.4097, 49650765224.4097, 
    49650765224.4097, 49650765224.4097, 49650765224.4097, 49650765224.4097, 
    49650765224.4097, 49650765224.4097, 49650765224.4097, 49650765224.4097, 
    49650765224.4097, 49650765224.4097, 49650765224.4097, 49650765224.4097, 
    49650765224.4097, 49650765224.4097, 49650765224.4097, 5903296507.56147, 
    43747468716.8482, 25642592941.4555, 8854944761.34219, 28715250851.106, 
    19860306089.7639, 2073933096.59516, 41794545276.1229, 49650765224.4097, 
    49650765224.4097, 49650765224.4097, 49650765224.4097, 49650765224.4097, 
    49650765224.4097, 49650765224.4097, 49650765224.4097, 49650765224.4097, 
    49650765224.4097, 49650765224.4097, 49650765224.4097, 49650765224.4097, 
    49650765224.4097, 49650765224.4097, 49650765224.4097, 49650765224.4097, 
    33938325327.8361, 20935514373.3036, 40795820463.0675, 34892523955.5061, 
    15274237177.4818, 4242843665.37253, 4242843665.37253, 4242843665.37253, 
    23554595083.7994, 4242843665.37253, 42750956463.7902, 28967627127.6403, 
    28967627127.6403, 48279378546.0671, 48279378546.0671, 48279378546.0671, 
    48279378546.0671, 48279378546.0671, 48279378546.0671, 48279378546.0671, 
    48279378546.0671, 48279378546.0671, 48279378546.0671, 48279378546.0671, 
    48279378546.0671, 48279378546.0671, 48279378546.0671, 48279378546.0671, 
    48279378546.0671, 48279378546.0671, 48279378546.0671, 48279378546.0671, 
    48279378546.0671, 48279378546.0671, 48279378546.0671, 48279378546.0671, 
    48279378546.0671, 48279378546.0671, 48279378546.0671, 48279378546.0671, 
    48279378546.0671, 48279378546.0671, 48279378546.0671, 48279378546.0671, 
    48279378546.0671, 48279378546.0671, 48279378546.0671, 48279378546.0671, 
    48279378546.0671, 48279378546.0671, 15377351998.8201, 15377351998.8201, 
    48279378546.0671, 13898719374.586, 5528422082.27687, 24609393423.8317, 
    23439205045.3634, 48279378546.0671, 48279378546.0671, 48279378546.0671, 
    48279378546.0671, 48279378546.0671, 48279378546.0671, 48279378546.0671, 
    48279378546.0671, 48279378546.0671, 48279378546.0671, 48279378546.0671, 
    48279378546.0671, 48279378546.0671, 48279378546.0671, 48279378546.0671, 
    48279378546.0671, 48279378546.0671, 48279378546.0671, 48279378546.0671, 
    13783329336.1499, 28967627127.6403, 48279378546.0671, 48279378546.0671, 
    48279378546.0671, 34479339689.2813, 2159999546.44369, 14419137616.7111, 
    11110100809.507, 34789442766.5701, 19578070893.07, 18739136709.5983, 
    46847841773.9957, 41688908497.6368, 41688908497.6368, 19687434907.517, 
    17527435361.0734, 36047844041.7777, 22157537531.2495, 12897333190.8973, 
    33267638340.7564, 46847841773.9957, 46847841773.9957, 46847841773.9957, 
    46847841773.9957, 46847841773.9957, 46847841773.9957, 46847841773.9957, 
    46847841773.9957, 46847841773.9957, 46847841773.9957, 46847841773.9957, 
    46847841773.9957, 46847841773.9957, 46847841773.9957, 46847841773.9957, 
    46847841773.9957, 46847841773.9957, 46847841773.9957, 46847841773.9957, 
    46847841773.9957, 46847841773.9957, 46847841773.9957, 46847841773.9957, 
    46847841773.9957, 46847841773.9957, 46847841773.9957, 46847841773.9957, 
    46847841773.9957, 46847841773.9957, 46847841773.9957, 46847841773.9957, 
    46847841773.9957, 46847841773.9957, 46847841773.9957, 41688908497.6368, 
    4319999092.8873, 10799997732.2181, 2159999546.44369, 28108705064.3974, 
    46847841773.9957, 46847841773.9957, 46847841773.9957, 46847841773.9957, 
    46847841773.9957, 46847841773.9957, 46847841773.9957, 46847841773.9957, 
    46847841773.9957, 46847841773.9957, 46847841773.9957, 46847841773.9957, 
    46847841773.9957, 46847841773.9957, 46847841773.9957, 46847841773.9957, 
    46847841773.9957, 46847841773.9957, 46847841773.9957, 39109441859.4573, 
    20370305149.8591, 28108705064.3974, 46847841773.9957, 46847841773.9957, 
    46847841773.9957, 45357938424.7518, 35766314628.4766, 19915447363.3629, 
    10946806485.9996, 40562126526.6142, 31593485649.251, 10946806485.9996, 
    33679900138.8638, 45357938424.7518, 45357938424.7518, 45357938424.7518, 
    22418951156.7134, 8757445188.7997, 40562126526.6142, 45357938424.7518, 
    45357938424.7518, 45357938424.7518, 45357938424.7518, 45357938424.7518, 
    45357938424.7518, 45357938424.7518, 45357938424.7518, 45357938424.7518, 
    45357938424.7518, 45357938424.7518, 45357938424.7518, 45357938424.7518, 
    45357938424.7518, 45357938424.7518, 45357938424.7518, 45357938424.7518, 
    45357938424.7518, 45357938424.7518, 45357938424.7518, 45357938424.7518, 
    45357938424.7518, 45357938424.7518, 45357938424.7518, 45357938424.7518, 
    45357938424.7518, 45357938424.7518, 45357938424.7518, 45357938424.7518, 
    45357938424.7518, 45357938424.7518, 45357938424.7518, 45357938424.7518, 
    45357938424.7518, 45357938424.7518, 38164220577.5454, 33368408679.4078, 
    4378722594.39982, 27631852358.5888, 27008869439.6768, 27214763054.8511, 
    45357938424.7518, 45357938424.7518, 45357938424.7518, 45357938424.7518, 
    45357938424.7518, 45357938424.7518, 45357938424.7518, 45357938424.7518, 
    45357938424.7518, 45357938424.7518, 45357938424.7518, 45357938424.7518, 
    45357938424.7518, 45357938424.7518, 45357938424.7518, 45357938424.7518, 
    45357938424.7518, 45357938424.7518, 45357938424.7518, 45357938424.7518, 
    40562126526.6142, 8757445188.7997, 4378722594.39981, 4378722594.39982, 
    7193717847.20638, 11989529745.344, 11989529745.344, 34305534094.4704, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 39371508497.9723, 
    11046107878.913, 28378408892.8697, 32711484146.3589, 41591516615.1768, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 32818425127.2787, 2209221575.78264, 
    8762304946.47628, 8762304946.47628, 26286914839.4287, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    43811524732.3812, 43811524732.3812, 43811524732.3812, 43811524732.3812, 
    41591516615.1768, 37151500380.7678, 34942278804.9852, 12999225760.4676, 
    21943053044.5177, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    25672467088.2849, 8442105467.1557, 8442105467.1557, 29764946328.4721, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 42210527335.7785, 
    42210527335.7785, 42210527335.7785, 42210527335.7785, 20976690174.4987, 
    6657944890.50751, 11096574817.5125, 25583463388.2483, 15273125701.0721, 
    40164287715.6849, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 16988975199.9031, 20580057747.2383, 2219396756.05894, 
    27156735899.2009, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 40556940878.3368, 40556940878.3368, 40556940878.3368, 
    40556940878.3368, 22880966619.5116, 6658190268.17683, 11865494955.4311, 
    36118147366.2189, 15538089618.9806, 40556940878.3368, 40556940878.3368, 
    32795148379.2897, 16261306989.6775, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 11196341026.5588, 10476164246.03, 10476164246.03, 
    12189052207.0223, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 30015851317.976, 
    34434338420.4239, 38852825522.8719, 38852825522.8719, 38852825522.8719, 
    38852825522.8719, 38852825522.8719, 38852825522.8719, 35427049600.8874, 
    32001273678.9029, 23311695313.7231, 18743084940.8361, 2209243551.22391, 
    26737471235.7076, 38852825522.8719, 6216666585.15317, 11448073662.9046, 
    34911650585.6817, 26157035388.7575, 26157035388.7575, 26157035388.7575, 
    34911650585.6817, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 34911650585.6817, 
    26157035388.7575, 15125314094.3679, 1554166646.28837, 22260182630.9477, 
    33991971092.3362, 4377307598.4622, 7354480862.92654, 8754615196.9243, 
    11731788461.3886, 33991971092.3362, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    7420060876.98264, 22260182630.9477, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 37100304384.9128, 37100304384.9128, 
    37100304384.9128, 37100304384.9128, 17882875032.4856, 32722996786.4507, 
    19151849338.3712, 22260182630.9477, 32722996786.4507, 19611455450.654, 
    10787241574.2492, 10787241574.2492, 4314896629.69962, 5605186972.50179, 
    23983530018.7909, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 30398697024.9032, 2157448314.84978, 
    21180936532.54, 35301560887.5667, 27596103538.6523, 2157448314.84978, 
    9106754092.03984, 17507835597.6902, 8629793259.39932, 16977046303.1636, 
    31097670658.1903, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    35301560887.5667, 33144112572.7169, 24514319313.3175, 7006483715.62725, 
    1401296743.12539, 4203890229.37632, 29642545453.1788, 35301560887.5667, 
    35301560887.5667, 35301560887.5667, 35301560887.5667, 35301560887.5667, 
    30986664257.867, 7006483715.62725, 1401296743.12539, 4203890229.37632, 
    15521921098.1521, 32498967401.3158, 9862905663.76422, 6346412250.57497, 
    10577353750.9583, 33458836041.2453, 33458836041.2453, 17614475916.8814, 
    7085633999.26671, 22881482290.287, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 33458836041.2453, 33458836041.2453, 28440160958.8267, 
    4230941500.38332, 7085633999.26671, 27112423790.6703, 33458836041.2453, 
    6691767208.24906, 4230941500.38332, 10455773520.063, 27185492188.222, 
    27185492188.222, 5437098437.64442, 2115470750.19167, 17220609125.8638, 
    30949498500.036, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    28021737603.6008, 6273343853.02326, 5018675082.41861, 2115470750.19167, 
    28882539583.1879, 33458836041.2453, 33458836041.2453, 33458836041.2453, 
    33458836041.2453, 31343365291.0536, 7085633999.26671, 15795848291.0203, 
    31343365291.0536, 4576296458.05741, 29345114173.0656, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 30459769912.354, 15600688173.1202, 
    6187764082.05668, 10312940136.7612, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    28230458433.7772, 26001146955.2003, 26001146955.2003, 26001146955.2003, 
    26001146955.2003, 26001146955.2003, 2229311478.57675, 21173966869.5622, 
    14565237239.7374, 10312940136.7612, 10312940136.7612, 4125176054.70443, 
    8250352109.40893, 10312940136.7612, 25092817070.0893, 27115802694.4888, 
    31574425651.6424, 31574425651.6424, 27115802694.4888, 8250352109.40893, 
    4125176054.70443, 10312940136.7612, 10312940136.7612, 27115802694.4888, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 31574425651.6424, 31574425651.6424, 
    31574425651.6424, 4458622957.15357, 6314885130.32842, 31574425651.6424, 
    31574425651.6424, 31574425651.6424, 15973737478.5221, 11848561423.8176, 
    10733905684.5292, 4125176054.70443, 8250352109.40893, 4458622957.15357, 
    4125176054.70443, 25653295999.3238, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 7893360401.06787, 17790406475.6704, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 21792782879.2684, 9993453650.31703, 27687452550.2728, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 26705840095.684, 
    12943285957.5549, 9993453650.31703, 9993453650.31703, 9826114432.83118, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 28669065004.8617, 26705840095.684, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    29650677459.4506, 29650677459.4506, 29650677459.4506, 29650677459.4506, 
    9993453650.31703, 1998690730.06342, 3931444761.82672, 19657223809.1336, 
    16707391501.8957, 4908062272.94438, 13858961713.8436, 5996072190.19022, 
    18842950572.0305, 26705840095.684, 28669065004.8617, 4948523037.30125, 
    1998690730.06342, 1998690730.06342, 1963224909.17776, 2567624564.9241, 
    15313091612.907, 23842601308.184, 27689988215.3633, 27689988215.3633, 
    18749630126.448, 6415011472.10356, 19160478520.0861, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 19995214401.005, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    18325742639.1675, 5771080360.76904, 20652184605.9817, 3847386907.17938, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 27689988215.3633, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 18749630126.448, 9618467267.94835, 15135325936.965, 
    20652184605.9817, 1923693453.58972, 1923693453.58972, 9618467267.94835, 
    9618467267.94835, 15135325936.965, 25978238505.414, 25978238505.414, 
    9364245576.19605, 13211632483.3754, 27689988215.3633, 27689988215.3633, 
    27689988215.3633, 18749630126.448, 7694773814.35869, 20652184605.9817, 
    9618467267.94835, 3847386907.17938, 855874854.974933, 855874854.974721, 
    4551013660.33228, 23486952350.4626, 25694800694.027, 25694800694.027, 
    16953347055.9581, 16959352576.0261, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 5212649718.3764, 8667532718.83779, 
    6946694887.43514, 21372433947.7118, 25419598734.7868, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 24219281921.8429, 
    11929423305.4286, 22006003763.5666, 24219281921.8427, 21879058614.0448, 
    2376892383.03431, 13245313292.9324, 21331663912.3518, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 20524079551.6815, 756384496.513565, 
    1749158312.19329, 8970354244.41275, 18271798157.9377, 25694800694.027, 
    25694800694.027, 25694800694.027, 20108534208.2463, 849649480.25639, 
    7970547523.02176, 23088716593.0081, 25694800694.027, 25694800694.027, 
    25694800694.027, 25694800694.027, 15152148517.4882, 10465135984.1837, 
    3933734759.27977, 7523017679.31969, 15531081895.7881, 16362326046.3087, 
    16432564018.795, 6578484479.92042, 4670098401.78983, 22339706625.9614, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    18952855988.0779, 1362653414.50392, 3427069789.23306, 3110717184.40749, 
    12288077714.7448, 22400559663.9041, 20815549552.2371, 22587421602.3663, 
    23375404988.385, 23649327120.6955, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 22295337156.8193, 14028676587.677, 2612753105.51673, 
    1225583342.78507, 3766873607.86844, 18335939960.7532, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23483339241.721, 19041563274.6126, 18861370200.9499, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23467712254.3051, 23577786617.0963, 8717199888.62121, 
    7833991541.1995, 4699700808.75031, 18392902360.3412, 23667600650.6443, 
    21805814880.5539, 13187553332.244, 679522255.264081, 7331093285.11295, 
    23654842447.0604, 23667600650.6443, 23667600650.6443, 23667600650.6443, 
    23667600650.6443, 23667600650.6443, 23667600650.6443, 20109261300.479, 
    5608143060.48052, 6821205606.23357, 12232791454.6109, 16869321775.1921, 
    21610913724.0339, 21592917995.0631, 20498982614.6496, 11168094858.8942, 
    8246205539.74249, 6361456011.5282, 1034687057.98075, 4710445.15715509, 
    2745697229.95101, 6887133.31899807, 1538019126.79614, 2477462816.76786, 
    3814314362.97885, 11694483564.2083, 12958383473.0687, 6559592538.60006, 
    18311298930.6103, 21470059675.9532, 16511650631.3304, 19883153925.9757, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 20789025685.1958, 21592917995.063, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 21595597604.1643, 21562943475.3861, 21610913724.0339, 
    20491885166.8398, 12903675952.6345, 13170473343.8549, 13347963200.3959, 
    4594901435.20991, 9015392832.88878, 13347963200.3962, 13170473343.8549, 
    5025814232.29711, 1630167110.03367, 5769623098.33847, 8520618372.5259, 
    16184269945.5707, 21463984809.3153, 21610913724.0339, 21592917995.063, 
    20498982614.6494, 18680719224.9201, 16730561405.3335, 14645224296.3858, 
    12422427833.037, 10058928156.4025, 8189993312.02375, 12180197899.7193, 
    13889237188.3308, 14441779152.4604, 15457094030.0056, 14261231504.1794, 
    12597640556.3107, 7891353948.76412, 10298387095.9138, 15865074661.3435, 
    14366981085.2655, 12139690128.9668, 13554441375.9423, 15171168736.891, 
    18455247294.3134, 20375176768.5054, 20630748303.2682, 21610913724.0339, 
    16818968511.5628, 7942994022.20166, 8734311362.06464, 20912241139.0084, 
    10555368449.0774, 8278544115.82541, 15864087402.1369, 21610913724.0339, 
    21556824054.9014, 18254473966.85, 764646842.881915, 12218352672.6424, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21610913724.0339, 21610913724.0339, 21610913724.0339, 21610913724.0339, 
    21587865958.9755, 13290104956.3094, 10043309207.3037, 6112051336.06095, 
    173511896.328593, 2139163512.55167, 594890272.571123, 4813121200.57235, 
    18558223402.3345, 4006990325.2342, 3916344234.84169, 16057512655.1958, 
    19318563019.1351, 3685297057.55917, 8241864280.73633, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 17750615091.6023, 
    392056952.660301, 6834950009.50953, 10960497179.6399, 12482862790.5513, 
    13872792027.6175, 15133159747.271, 16268225313.1675, 16594352243.7529, 
    7964407567.30501, 122397177.9736, 667425229.862553, 955591455.117576, 
    2234115697.98869, 5918901779.65834, 3117171773.38077, 2139163512.55946, 
    594890272.571113, 776664092.989111, 9517145621.53167, 12415118165.9307, 
    10322247363.8497, 19438114723.9258, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19194324309.4753, 3738793965.39504, 942132079.820964, 
    7489201830.7119, 15748926769.6277, 15121343377.2022, 871441353.651519, 
    13085220828.2727, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19228902971.5441, 12412873656.8389, 5330902247.16945, 
    111788325.441386, 1054098190.7576, 17838878447.5, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19527302289.9998, 19527302289.9998, 
    19527302289.9998, 19527302289.9998, 19197714480.7758, 6567503859.49613, 
    538525803.71136, 11204183255.0186, 13502136933.4364, 1508915725.52588, 
    2229524623.649, 5109809674.25509, 71625395.7381112, 449431133.320748, 
    1489032083.37468, 12298054479.4126, 11718637446.5849, 12367369471.8185, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 13877928980.2487, 11331224160.5156, 
    6993276250.19654, 2949543688.32432, 5559729768.29254, 8018726080.42385, 
    2934331879.25452, 1506370619.05243, 6174373140.1154, 4870380867.3698, 
    3702999539.4386, 2667399985.45729, 598381498.84628, 444103701.478904, 
    11049184794.3143, 14127834115.424, 11078480495.3158, 9920948777.19226, 
    3424356448.26897, 3488666850.21017, 5796244477.83205, 7767340043.75177, 
    1791796495.88034, 1113432615.29749, 12298054479.4124, 12277208215.6665, 
    13711154286.7809, 4626290523.04475, 1623757012.8143, 7922014819.08065, 
    9091869980.9416, 8617548800.07451, 6820771883.05755, 2076648695.53807, 
    6698774073.04278, 17374232424.7742, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 17419362268.9296, 17419362268.9296, 
    17419362268.9296, 17419362268.9296, 10005124093.8306, 15914383.7275346, 
    2775552891.106, 9401477771.27636, 8049929997.3472, 6992277446.12201, 
    4973223170.54911, 126553906.525535, 46415086.5523994, 7090117628.32968, 
    8875935041.10666, 12279066153.8603, 13086831685.2862, 12828210240.3574, 
    15118515953.2275, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    14420604374.0182, 5483756119.24378, 51822629.5140081, 640115627.532849, 
    7608757323.2762, 9246384036.81436, 10372059135.1033, 4837991613.5002, 
    5176789279.88169, 930662031.230483, 417075478.271312, 6129858745.72945, 
    6324968997.50866, 9468783921.48417, 8723310854.67286, 9762660834.99837, 
    11349613816.6761, 10277503167.9502, 6316917206.02679, 6386704279.17343, 
    13093129059.3211, 3658395586.21854, 3221689419.30748, 10690391486.0232, 
    15072601047.0027, 13326711869.0605, 13748541502.0964, 12478527673.065, 
    1145189957.39974, 1808130373.88102, 2024205293.62305, 4580762095.69292, 
    5187219478.12986, 8978019688.93456, 14828334317.1595, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    15289719891.5999, 15289719891.5999, 15289719891.5999, 15289719891.5999, 
    10276198021.7206, 4418821677.75221, 859949263.074625, 7598690407.25748, 
    10885599222.7918, 7333717261.21515, 6591131069.00275, 2720995424.46681, 
    50977672.1746417, 706855736.218169, 103838582.715547, 66846344.6646293, 
    2402107067.79995, 5331209189.57717, 4593754600.39129, 4538789156.51487, 
    1160867855.56029, 895904772.221222, 4694017319.28048, 4158156933.67979, 
    229984186.987567, 2123633631.31493, 4291765471.25796, 4291765471.25796, 
    5952764573.13931, 6212540814.2187, 5996713187.84684, 10092634917.327, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 9767398175.37204, 
    1478117095.79851, 826412938.04413, 9077104919.55163, 12994606455.0839, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 13141028427.2218, 13141028427.2218, 
    13141028427.2218, 13141028427.2218, 5230007080.50411, 1013138432.4626, 
    8087609624.64994, 7572547211.59138, 6703075023.87572, 6351442695.58753, 
    8513436297.27524, 3432460258.43351, 41810879.4074752, 1444554249.11809, 
    3146312860.00849, 1750656533.82562, 1541222179.18314, 3094720547.55575, 
    2905936038.84418, 2665039479.94633, 883983261.389403, 191806505.092574, 
    5269186194.44947, 8627483873.4555, 9954664514.97536, 7828250510.23732, 
    5778750279.48653, 2788031449.23336, 611889535.478295, 2518707669.68707, 
    3581544054.19524, 5011306624.78963, 5071892667.35915, 10657380130.2225, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10920377367.1557, 8087285125.3005, 3869454895.18043, 
    298503060.881661, 740480057.471925, 6175959643.10779, 10742615937.0253, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    10975964877.7963, 10975964877.7963, 10975964877.7963, 10975964877.7963, 
    8595542346.16688, 2797872551.98662, 131614991.8018, 1225570182.58736, 
    2364821153.62565, 589670242.589798, 103085954.921991, 93034863.9796758, 
    1054987094.45796, 2587701086.98983, 1864297442.59602, 32043176.6406526, 
    3004453836.81918, 4511053605.69711, 4190484509.76999, 6325759004.06176, 
    8787246866.57545, 8797226642.9036, 8589874130.6553, 8097264479.69153, 
    4989141722.20048, 2607678092.87671, 699108410.087622, 1023677.07039754, 
    986479475.635109, 2656667517.22495, 4096506130.04143, 5342331534.61792, 
    6423498484.53633, 7363443596.42065, 8182553501.70449, 8756114186.16336, 
    8797226642.9036, 8797226642.9036, 8797226642.9036, 8797226642.9036, 
    8797226642.9036, 8797226642.9036, 8695384737.31328, 8420069132.42867, 
    7047209334.48159, 4724298397.75764, 4717944377.39766, 3074024056.79447, 
    559350932.776624, 269675403.267611, 1153050.7646866, 491068003.467734, 
    2166183028.60623, 1969352673.52792, 1279779249.71046, 142226953.325068, 
    141393683.628623, 723474919.522283, 1267076982.4447, 1740669545.31719, 
    2150481113.61707, 2504513530.46523, 2807953527.99078, 1167652719.74651 ;

 tile1_distance =
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000841027571416003, -0.00647256284921793,
  2.02680978575187e-16, -0.0103889353725783,
  -1.51996163746982e-16, -0.0103889353725777,
  2.02680978575187e-16, -0.0103889353725783,
  -1.51996163746982e-16, -0.0103889353725777,
  2.02680978575187e-16, -0.0103889353725783,
  -2.02661551662642e-16, -0.0103889353725777,
  1.52015590659526e-16, -0.0103889353725783,
  -2.02661551662642e-16, -0.0103889353725777,
  1.52015590659526e-16, -0.0103889353725783,
  -1.51996163746982e-16, -0.0103889353725777,
  2.02680978575187e-16, -0.0103889353725783,
  -1.51996163746982e-16, -0.0103889353725777,
  2.02680978575187e-16, -0.0103889353725783,
  -2.02661551662642e-16, -0.0103889353725777,
  1.52015590659526e-16, -0.0103889353725783,
  0.00046904711303759, -0.00225077484656944,
  8.70305234902186e-21, -0.00133932228146305,
  2.2680154421551e-17, -0.00133932228146305,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -9.65457151894165e-05, -0.000777390578489801,
  0, -0.00133932228146305,
  -0.000935856603785424, -0.00497643624457078,
  -1.51996163746982e-16, -0.0103889353725777,
  3.5463828849708e-16, -0.0103889353725783,
  -1.51996163746982e-16, -0.0103889353725777,
  3.5463828849708e-16, -0.0103889353725783,
  -1.51996163746982e-16, -0.0103889353725777,
  0.000747259341699632, -0.007147621063059,
  0, -0.00133932228146305,
  6.5430558101785e-05, -0.00105369977971459,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.003802572397468, 0.00237538176162855,
  -8.86452399801261e-17, -0.0105324026284572,
  -8.90879553545946e-17, -0.010532402628457,
  1.36220115221093e-19, -0.0105324026284572,
  0.00109252041556442, -0.00513419425036288,
  5.92270150459521e-17, -0.00153437536304701,
  -5.92270150459521e-17, -0.00153437536304701,
  0.000125269156276316, -0.00057989605621156,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000127615555379234, -0.000886137012599431,
  -0.000873957280668704, -0.00729369643538091,
  -0.00307296182761978, -0.0105324026285623,
  0.00409728243682734, -0.0105324026287401,
  -8.91220103833998e-17, -0.010532402628457,
  9.86965519132316e-17, -0.00153437536304701,
  8.20049888897309e-05, -0.00028471315921097,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000662784075248795, 0.00201400286467868,
  -0.000993955532337538, 0.00735999536815024,
  6.32996910425545e-16, 0.0156276438892191,
  0.00234496877735149, -0.0106884896865793,
  3.98409441571039e-17, -0.0106884896865955,
  0.00100524854562919, -0.00744361734398002,
  -3.70642879100138e-17, -0.00172945690614368,
  -1.07196555338738e-16, -0.00172945690614368,
  -3.70642879100138e-17, -0.00172945690614368,
  -1.07196555338738e-16, -0.00172945690614368,
  -1.75397922376403e-17, -0.00172945690614368,
  3.70642879100138e-17, -0.00172945690614368,
  1.07196555338738e-16, -0.00172945690614368,
  -0.000625071921552112, -0.0026177350490133,
  -9.01521835742872e-17, -0.0106884896865955,
  0.00100524854562933, -0.00744361734398002,
  0.000104323491002423, -0.000317759143315,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -7.21169708634574e-17, -0.00172945690614368,
  -3.70642879100138e-17, -0.00172945690614368,
  -7.21169708634574e-17, -0.00172945690614368,
  -3.70642879100138e-17, -0.00172945690614368,
  0.000159733112991046, -0.000648708571839629,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00351745316602714, -0.0106884896865589,
  0.0011724843886758, -0.0106884896865898,
  0.00107285632305542, -0.0037622786009508,
  0.000104323491002423, -0.000317759143315,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00020306152432128, -0.00110000188880299,
  1.58394890474117e-17, -0.00192454349003279,
  -0.00415439729867557, 0.0049568574612231,
  0.0013192182159598, -0.0108530285837203,
  -4.21325723614263e-17, -0.010853028583717,
  2.85162457445051e-16, -0.0108530285837161,
  -2.85385714627729e-16, -0.010853028583717,
  4.1909315178748e-17, -0.0108530285837161,
  0.00263843643191924, -0.0108530285837276,
  0.000895393442020853, -0.00183026463659575,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.0013192182159598, -0.0108530285837203,
  -4.21325723614263e-17, -0.010853028583717,
  0.000705304704323412, -0.00280075081585096,
  -2.79450598097878e-17, -0.00192454349003279,
  2.79450598097878e-17, -0.00192454349003279,
  0, 0,
  0, 0,
  1.34672373891069e-16, -0.0110235014048152,
  6.74396219485232e-17, -0.0110235014048148,
  -3.39783984817329e-17, -0.0110235014048152,
  6.78533619604773e-17, -0.0110235014048148,
  -6.76982094559945e-17, -0.0110235014048152,
  6.78533619604773e-17, -0.0110235014048148,
  -3.2279106937658e-17, -0.0110235014048152,
  3.56259725243137e-17, -0.0110235014048148,
  -3.2279106937658e-17, -0.0110235014048152,
  3.56259725243137e-17, -0.0110235014048148,
  -3.2279106937658e-17, -0.0110235014048152,
  0.00158975698599842, -0.00560959476647871,
  -1.45134583707892e-17, -0.00211962057082271,
  0.000156737325602864, -0.000381658445970601,
  -1.45134583707892e-17, -0.00211962057082271,
  4.34736976619657e-17, -0.00211962057082271,
  0.000241115863002936, -0.000782829107817795,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000786970441461855, -0.00298343389500833,
  -6.7025881936569e-17, -0.0110235014048148,
  0.00135486901112635, -0.00410250555637748,
  0.000156737325602864, -0.000381658445970601,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -7.24783885867434e-17, -0.00211962057082271,
  7.24561627699428e-17, -0.00211962057082271,
  -2.06870005977065e-19, -0.0110235014048152,
  6.74396219485232e-17, -0.0110235014048148,
  -0.00439301081016628, -0.0110235014047964,
  0.00439301081016624, -0.0110235014047959,
  0.00128211246787687, -0.00774883241669322,
  4.86668374474119e-17, -0.00211962057082271,
  0.000241115863002997, -0.000782829107817795,
  0, 0,
  0, 0,
  0, 0,
  6.88803259851298e-17, -0.0110235014048152,
  -3.16067794182295e-17, -0.0110235014048148,
  0.00160765899562398, -0.0111982975267613,
  0.00321531799124775, -0.0111982975267604,
  1.58565511505501e-16, -0.0111982975267626,
  0.00150048752085241, -0.00427174532432906,
  2.67578813540139e-17, -0.00231467869401381,
  0, 0,
  0, 0,
  -0.000186737510290506, -0.00041249829650547,
  -1.34405947815093e-17, -0.00231467869401381,
  -4.01573733991882e-17, -0.00231467869401381,
  -0.00150048752085238, -0.00427174532432906,
  -3.21010301579943e-17, -0.0111982975267635,
  1.58177583648606e-16, -0.0111982975267626,
  0.00160765899562402, -0.0111982975267613,
  0.00150048752085238, -0.00427174532432906,
  2.67578813540139e-17, -0.00231467869401381,
  0, 0,
  -0.00028794937894355, -0.000848096904289219,
  -2.67578813540139e-17, -0.00231467869401381,
  0.000296244367257466, -0.00130879218270574,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000186737510290506, -0.00041249829650547,
  -4.11027363348907e-20, -0.00231467869401381,
  -6.95405847678311e-18, -0.00231467869401381,
  2.67578813540139e-17, -0.00231467869401381,
  -0.000186737510290506, -0.00041249829650547,
  2.67578813540139e-17, -0.00231467869401381,
  0, 0,
  0, 0,
  0, 0,
  -0.000203354293550835, -0.00179681735172132,
  -2.67578813540139e-17, -0.00231467869401381,
  6.95405847678311e-18, -0.00231467869401381,
  -0.00176475933745515, -0.0057673081513141,
  -9.4363451189512e-17, -0.0111982975267626,
  3.1325174444206e-17, -0.0111982975267635,
  -3.13251744442059e-17, -0.0111982975267626,
  0.00328715439556407, -0.00231467869401336,
  0.000296244367257475, -0.00130879218270574,
  0, 0,
  0, 0,
  3.52797269557491e-17, -0.0113763388323844,
  1.19580475144781e-16, -0.0113763388323844,
  -0.00174900597690388, -0.0113763388323807,
  -8.98231218829461e-17, -0.0113763388323844,
  -0.00349801195380749, -0.0113763388323747,
  0.00524701793071145, -0.0113763388323624,
  -1.25006221349597e-17, -0.00250971147676093,
  1.25006221349597e-17, -0.00250971147676093,
  -1.25006221349597e-17, -0.00250971147676093,
  -0.00157915761507213, -0.00805554410828924,
  -5.98820812552974e-17, -0.0113763388323844,
  1.19580475144781e-16, -0.0113763388323844,
  -1.19580475144781e-16, -0.0113763388323844,
  5.95147065236698e-17, -0.0113763388323844,
  -0.00174900597690369, -0.0113763388323807,
  -0.00174900597690384, -0.0113763388323807,
  -8.96394345171323e-17, -0.0113763388323844,
  8.96394345171323e-17, -0.0113763388323844,
  2.99410406276487e-17, -0.0113763388323844,
  -0.00699602390761477, -0.0113763388323256,
  0.00524701793071078, -0.0113763388323624,
  0.00188778160718909, -0.00218986953459233,
  0, 0,
  -3.17265386929203e-17, 0.0149720637764361,
  -0.00741489283440082, 0.0149720637765796,
  0.00377640492436723, -0.0115568764838534,
  4.53196279150453e-17, -0.0115568764838549,
  0.00180092245015882, -0.00460804381674307,
  -0.0076915568602264, -0.00270471446921161,
  0.0100598624068692, 0.0140713850258246,
  -2.39139513053582e-17, 0.0140713850257925,
  -1.80962443210508e-16, 0.0140713850257927,
  -0.00502993120343444, 0.0140713850257976,
  0.00378991243458344, 0.0046592334222626,
  0, 0,
  -0.00218289951798814, -0.00245068912220681,
  -0.00509200918354315, -0.0124823876706783,
  0.00827666594417081, 0.013700451790552,
  0, 0,
  0, 0,
  -0.00813655246754144, -2.22044604925031e-16,
  0.008148921039913, 0.00117571017422036,
  -0.00271630701330447, 0.00117571017422113,
  0.00850144301375317, 0.00079039807666903,
  0.00849324022692447, 1.4432899320127e-15,
  0, 0,
  0, 0,
  -0.00276538929388932, 0.00275881786357524,
  -0.011503301136772, 0.0135136099914021,
  0.00298921849691848, 0.0133260244548715,
  0.00871306733904991, -0.0130480411670464,
  0, 0,
  0, 0,
  0, 0,
  -0.00739025861552715, 0.000201195719833125,
  0.0122333407211158, 1.81991816727844e-05,
  0.00137569652936377, 2.00238266268027e-06,
  -0.00921626134475611, 0.00446276028894699,
  0, 0,
  0, 0,
  0, 0,
  -0.00451570512760892, 0.00661272685561609,
  0.00135443335269903, 0.00725001390666069,
  -0.0128192814076929, 0.0129490055497028,
  0.0031256148063672, -0.0134275349928427,
  0.000148567515104016, 0.000767558637041921,
  -0.00880987128708944, 0.00783511380293145,
  0.00415491699688499, -0.00186100178411819,
  0, 0,
  0, 0,
  0, 0,
  -1.63046970171339e-17, -0.00484723462230119,
  -0.013024217981644, -0.00484723462230086,
  0.00921608622696648, -0.00825754653853505,
  -0.00319146487794225, -0.00128923663372871,
  -0.00330676335836679, 0.0127597237979629,
  0.00654002951523204, 1.11022302462516e-16,
  0, 0,
  0, 0,
  0, 0,
  -7.45685607731083e-17, 0.0127597237979628,
  -0.0132270534334662, 0.012759723797962,
  0.00340463199710865, 0.0125700079533879,
  -0.0034046319971087, 0.0125700079533883,
  0.010067910581089, -0.00504175533107409,
  -0.00223527555311485, 0.000839527155031772,
  -0.0136185279884344, 0.0125700079533967,
  0.00673980141445895, 5.55111512312578e-16,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00446648270588346, 0.00671010518384474,
  -0.00340463199710872, 0.0125700079533883,
  -1.39202488753246e-17, 0.00369560432081484,
  0.000597779069415395, 0.000610243832200541,
  -0.00059777906941539, 0.000610243832200541,
  1.39202488753246e-17, 0.00369560432081484,
  0.0104949170722946, 0.0123799068809152,
  -0.00504825639071548, -0.00793814970460927,
  -0.0137132575335287, -0.0139992034806229,
  0.00777955530398675, -0.00305947341796198,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000597779069415386, 0.000610243832200541,
  -0.0139017242803413, 0.00369560432081806,
  0.00717533806362134, 0.0121894621555841,
  -0.00717533806362113, 0.0121894621555845,
  0.00344818163487326, 0.00876576126330852,
  6.77195592185708e-18, 0.00350296830735197,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0107630070954318, 0.0121894621555656,
  0.00472294018180723, -0.00396789428775068,
  0.0141731435512379, -0.00543065996801262,
  0.00094270822402566, -0.000800736224458531,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00439122695462554, 0.00673026709890101,
  -0.010763007095432, 0.0121894621555656,
  0.00365189814417321, 0.003310052279205,
  -6.92259778820377e-18, 0.00331005227920345,
  6.2005480290863e-18, 0.00331005227920345,
  -0.00201236971890476, 0.00408668687050695,
  -0.0073452238496415, 0.0119987093638553,
  0.00728782031798936, 3.10862446895044e-15,
  -0.000875879669139759, 0.00116336457360822,
  -4.9123960422786e-18, 0.00331005227920345,
  -0.00350289616802813, 0.00511255096737739,
  -0.0110178357744622, 0.0119987093638676,
  0.0110178357744622, 0.0119987093638678,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00739821193900336, 0.00290308600021394,
  0.00364391015899449, 1.11022302462516e-15,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00284852831690171, 0.00233491083992199,
  -0.0146904476992832, 0.0119987093639058,
  0.015012118888663, 0.0118076791352705,
  0.0022976594459775, 0.000900242321607125,
  0, 0,
  0, 0,
  0, 0,
  -0.000840044194991332, 0.00110495364304974,
  -0.0112590891664971, 0.0118076791353009,
  0.00407722517072194, 0.00212998821319776,
  0, 0,
  0, 0,
  0, 0,
  -0.000873146224592913, 0.00172274168585096,
  0, 0.00311687794791271,
  6.21639461346925e-18, 0.00311687794791271,
  0.000873146224592913, 0.00172274168585085,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000539573576337367, 0.000532296805711652,
  -0.0149337442958426, 0.00311687794789328,
  0.00372631727830079, -1.11022302462516e-15,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00411815355878268, 0.00390936779992823,
  0.0105953664187832, 0.00471132433195931,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00753276722959315, 0.00295527613274682,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0152163347363459, 5.77315972805081e-15,
  0.00537552315420169, -0.00239027439282158,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0114864309470561, 0.0116101901586175,
  0.000748419816704014, 0.000972340250275872,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00048327607599959, 0.000470900927061813,
  -0.015530176480574, 0.00269279643967801,
  0.0116476323604304, 0.00269279643968007,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.015508449519868, -3.27515792264421e-15,
  0.0116313371399012, -1.16573417585641e-15,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00451356590219111, 0.00123545544316694,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00371905788522579, 0.00654613277119059,
  0.0118956763909707, 0.010716381606046,
  -0.00693993841778243, 0.00488986226211685,
  0.0118359368599039, 1.88737914186277e-15,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00135088643164372, -0.000912723289041073,
  -0.0157298012656, -0.00692173735436924,
  0.0118359368599041, 1.88737914186277e-15,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00217577624857944, 0.000957427972564318,
  -0.0158609018546282, 0.0107163816060539,
  0.0120334525281658, 0.0014648402341178,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.00702759631000854, 0.00300976351499871,
  -0.000268172291474939, 0.000273229515340534,
  -0.0160446033708879, 0.00146484023412674,
  0.0120257950600073, 4.9960036108132e-15,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0108015192320728, -0.00124075498709747,
  0.0119409966010901, -0.0162215750480632,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000282444423375918, 0.0011510831709749,
  5.5997344208541e-18, 0.00966543883719972,
  -0.0161009129700272, 0.00966543883722959,
  0.00645160441477291, 0.00283063465503436,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.00712532107552869, -0.00300937554608172,
  0, 0,
  -0.0141315039044774, 0.00276185949977864,
  -0.0122300907723128, 0.00614557131775512,
  0.0121161858800779, -0.0175593638723587,
  0.00299551044031185, -0.00383834134349675,
  0.000557896532467144, -0.00107334510099755,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0033803931226346, -0.00327466044855063,
  -0.0121161858800817, -0.0175593638723633,
  0.00405185402782281, -0.00950653280283514,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00679490105831814, 0.00112789385022627,
  0.0165132341782858, 0.00566928616002543,
  0.00112584715992544, 0.000822715837849708,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00779174984370804, 0.00771329459413317,
  0.0123603585756141, 4.44089209850063e-16,
  0, 0,
  -0.00824023905040938, 2.22044604925031e-16,
  0.0123083906711995, -0.0119925194159946,
  0.00469843211537228, -0.00465112352980157,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00352182766115464, -0.00280611159565131,
  -0.0164111875615991, -0.0119925194159911,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.0166728622945793, 8.93729534823251e-15,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00201806386807772, 0.000982698576508512,
  2.06893314198155e-17, 0.00954761275910132,
  0.0124733667980866, -0.00809856086362482,
  0.000374483065655363, -0.000487127442375779,
  -0.000770351988651717, 0.000934454392040263,
  0.0166311557307828, -0.00809856086361482,
  0.00317722675887285, -0.00362813945402962,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000245990213456858, -0.000239987988484236,
  -0.0020900725790464, -0.00605123404274166,
  0.00276971691097861, -0.00282639737142337,
  0, 0,
  -0.0125046467209344, 3.38618022510673e-15,
  0.0166448721121761, -0.00551897463434453,
  0.00266415527062697, 0.00360846193586067,
  0.0137179436210933, 0.0111773672371085,
  0.00319909495823622, 0.00568660832534701,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0125147432236343, 0.00257524023494959,
  0.0168444793595266, -1.46549439250521e-14,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.0108227238091771, -0.00891518319080159,
  0.00119800593907348, -0.000836613200063174,
  0.0125908223158657, -0.0123149913376774,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00872297614880497, -0.00286128806405656,
  0.0168444793595264, -1.46549439250521e-14,
  0, 0,
  -0.0125908223158656, -0.0123149913376774,
  0.0126518218266421, 0.00534504223463717,
  0.00173427147880127, 0.0016962782654516,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0126333595196449, -5.44009282066327e-15,
  0.0169252950128165, -0.0171820213876355,
  0.00410294929386811, -0.000118335576312856,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.00690390039811719, -0.00700888904713193,
  7.19579352490323e-17, -0.0171820213875951,
  -1.51911196636847e-16, -0.0171820213875966,
  0, 0,
  0, 0,
  -0.00622067968847633, 0.00255529498762005,
  0.0169951153252319, -1.19348975147204e-15,
  -0.0089736322791487, -0.00322379698432823,
  0.00622067968847644, 0.00255529498762,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00903540398540835, 0.00277445913183752,
  0.00428114559636813, 2.77555756156289e-17,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00429176369832629, 0.0127869540902144,
  -0.00885080647892614, -0.0118053464404634,
  7.72752798023781e-17, -0.0166104622237646,
  -0.0042667958708871, -0.0166104622237638,
  0.0171245823854724, 7.49400541621981e-16,
  -0.0171245823854733, 7.49400541621981e-16,
  -0.0128752910949784, 0.0127869540902144,
  0.0171481109048239, 0.00694397278647102,
  0.00145913973717534, 0.000914447586569417,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000206651971111824, 0.000201121922836806,
  -0.0123893489004502, 0.00538725803945972,
  0.00430817978254438, 2.77555756156289e-17,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00423045650931243, -0.00221638386578282,
  0.00863340876103138, 0.012547192076286,
  0.00403207889688171, 0.009160390865808,
  -0.00431670438051591, 0.012547192076286,
  0.0115754536838799, -0.00509477371678058,
  -0.0129286140381685, 0.00168762141953729,
  0.0101013647400792, 0.00374165434428791,
  -0.0172327191301782, 5.55111512312578e-17,
  0.012333584912331, 0.00536822004101878,
  -0.00461559712811289, -0.00376746411613021,
  -0.0128888664429719, -0.0166854484592409,
  0.0101013647400791, 0.00374165434428791,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00234137677012048, 0.0019733840245196,
  0.0173441042097491, 0.011670002155229,
  0.00263826309560813, 0.000910807402032782,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00865969537244044, 1.47104550762833e-15,
  0.00916150324949214, 0.00359883558043586,
  -0.00194013630446724, -0.00169759479106453,
  8.68377746458004e-18, -0.00535937034208663,
  -0.00865408113459215, -0.00535937034208429,
  0.00864055754162988, -0.0170462054994333,
  7.02979268406852e-18, -0.0170462054994755,
  -0.00432027877081515, -0.0170462054994599,
  0.0043239738867626, -0.0108291274826098,
  0.0130157213204182, 0.0169736796121993,
  0.00433019298636646, 0.000615122718007788,
  0.000183115178355478, 0.000240834687290581,
  -0.000123826245597522, 0.000488572090058301,
  -0.00248344906844709, 0.000915717878000211,
  -0.011779298761685, 0.00972251565471263,
  -0.0130157213204182, 0.0169736796121989,
  -0.0130071225419589, 0.0110068898372211,
  0.0130157213204182, 0.0169736796121993,
  0.000183115178355486, 0.000240834687290581,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.0136264188089776, 0.00405681182720323,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00610468856198326, 0.00167408096109334,
  0.0174052724367842, 0.0140692209970093,
  0.0045133698309543, 0.00694200728608836,
  -0.0130383668830338, -5.55111512312578e-16,
  0.0130436737280017, 0.00445376961272437,
  0.00362353535453495, 0.0123458138551645,
  -0.0173988397915046, 0.00936889921267522,
  0.0130365858485129, -0.00105494665641123,
  -2.54193035757269e-18, 0.00936889921267843,
  0.00206350573567965, 0.000983473983302049,
  0, 0,
  -0.0011511176376752, -0.00124064540380614,
  -0.00743331819810547, -0.00986452301740963,
  0.0130226387631823, -0.0131998245068008,
  -0.00390883872502863, -0.0082794635414684,
  0.0130383668830338, -5.68989300120393e-16,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00180151107745788, -0.000970074781852404,
  -1.77193295980234e-18, -0.00827946354146736,
  0.0130813180586132, 0.0165888597113438,
  0.00172668442283236, 0.00165227140274775,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0130813180586133, 0.0165888597113438,
  0.0129094811497179, 0.00448916763256778,
  0, 0,
  -0.00621601652542828, 0.00161134759287272,
  0.00151163391969666, 0.00809182728293253,
  3.05433644883269e-18, 0.00515232718864796,
  -0.0130716394205585, 0.000905145496472068,
  0.0130709499535103, -4.02455846426619e-16,
  -0.00408150043753999, -0.000211967582318742,
  -0.0174109224479353, -0.0167491001703783,
  0.00435422676437261, -0.0115933887468934,
  0.00435727760643271, 0.000490142350745779,
  0.00509346989580011, -0.00162349760743991,
  0.000883820570706858, 0.000753690500485092,
  0.000320713552997988, -0.000406707650893845,
  -0.000320713552997986, -0.000406707650893845,
  -0.00239142769425058, -0.0053700903986261,
  -0.0140198426988652, -0.0136038797554711,
  0.0130760146822948, 0.00815197616136229,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000792809657242775, -0.00164587297527988,
  7.50468637909005e-19, -0.0046630297322219,
  -0.0104600586469341, -0.0131339678137549,
  0.0130872516500458, 5.58580959264532e-16,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00491640671745635, 0.00286325072872732,
  -0.0174531934586843, 0.0147297407813946,
  0.00191212028103288, 0.00175712501109269,
  -0.00330561037504302, -0.00221046207102306,
  -0.0130828596186457, -0.0152845650227574,
  0.0130887082689936, 0.00562611620065432,
  0, 0,
  0, 0,
  -0.00498907857663337, 0.00109799834686511,
  0.0130841387164986, -0.0120235466436983,
  -0.00387489091353532, -0.00215094515417618,
  -0.00173754653099382, -0.00508852182857778,
  0.0174507011085068, 0.00412484482448047,
  -0.0174507011085068, 0.00412484482448043,
  0.0114936930506627, -0.00170190747430914,
  -0.00939749172092263, -0.00473545806307799,
  0.00872190641243054, -0.0152845650227598,
  -0.00872190641243048, -0.0152845650227598,
  0.0130860465084483, -0.00587200439000862,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000927114657252312, -0.00104325958900872,
  -0.00119349755768086, -0.00452887489094169,
  -0.00313109762331397, -0.00991022843348854,
  0.0130887082675291, -0.00562610922035122,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00759368292481682, 0.00458539271727791,
  0.0174503886225849, 0.000245510702510675,
  0.00296582857588982, 0.00381623503435758,
  0, 0,
  -0.0100451177721033, -7.43067534797366e-05,
  0.0130872516500458, -5.55111512312578e-16,
  0, 0,
  0, 0,
  -0.00124418765291922, 0.000839517521394339,
  -0.0174480620088773, 0.00587201137230006,
  -0.00187649544090182, -0.00878793373597745,
  0.00395373752651506, -0.00356653888121045,
  0.0174505753449234, -0.00236595337012652,
  -0.00951268901618319, 0.00263016755466915,
  0.00479635525319509, -0.00351277379116736,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00178050173762006, 0.000175785922105497,
  0.0130581918296153, 0.0167491071519647,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00840509331544479, 0.0040313113650696,
  -0.0174109224394868, 0.0167491071519777,
  0.0158249822495276, 0.00614141422044687,
  -0.000634846210203235, -0.00137881313328618,
  0.00172668177383135, -0.00165226979172139,
  -0.00976740212433143, -0.00301992344031832,
  0.0130813180552598, -0.0165888527301445,
  0.0070793701654635, -0.0146968289993651,
  0.00318762589251227, -0.00123706495698083,
  0, 0,
  -0.0174279332713477, 1.00613961606655e-15,
  -0.00436043935175337, -0.0165888527301445,
  0.017432911808227, -0.00515232021047848,
  0.00107975361564088, -0.000774915929210286,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00886831005231726, -0.000592748112752582,
  -0.0130226387540606, 0.0131998314901759,
  0.00201346398240683, 0.00502072486418279,
  0.00120421495533712, 0.00194680755495411,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0106684850168405, 0.0042636812649321,
  0.00293534604285352, -0.0035393621479598,
  -0.0173988397815741, -0.00936889223455997,
  0.0030143849354644, 0.0021642399124235,
  -0.0173844891773788, 1.4432899320127e-15,
  0.0130491298361806, -0.00936889223456192,
  0.00146167884147311, -0.00148156719729164,
  -0.0105840938265793, -0.000459143956748426,
  -0.0130226387540605, 0.0131998314901759,
  0.00434612229434476, 8.32667268468867e-17,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0014616788414731, -0.00148156719729164,
  -0.0013992811886928, -0.00512019845762295,
  -0.0173988397815748, -0.00936889223455997,
  0.00158729588096676, 0.00699496938533839,
  -0.00158729588096676, 0.00699496938533839,
  -1.77226289770592e-18, 0.0082794705268015,
  -0.00346288478397193, 0.00946329658056315,
  -0.000200449220343439, 0.000392105750117513,
  -1.13072565727916e-18, 0.000663731409923651,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00455163690748776, 0.00217360381813118,
  0.0172811150662107, 0.0170462124809187,
  -0.0172811150662104, 0.0170462124809149,
  -0.0044889101114772, 0.000361824813403105,
  0.0114126683138639, 0.0119496209670181,
  -0.00812288209536209, -0.00367813529267226,
  -0.0173542950809055, -0.0169736726312004,
  0.00895743015636026, -0.0107180941843344,
  -0.0173382296632994, -0.00899184580064846,
  0.0172958955144068, 0.0108291414450983,
  0.00559558358273833, 0.00433228420394076,
  -0.00882380634315976, 0.00260555681891587,
  0.0172811150662094, 0.0170462124809187,
  0.0101755645756484, 0.0121693554067356,
  0.0135438482319826, 0.00790112677145947,
  0.00125992374354373, 0.000847740756430598,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00552129659076203, -0.0044268418347258,
  -0.0149790482662629, -0.0126344690125169,
  0.0172811150662112, 0.0170462124809187,
  0.00568936712019418, 0.00297790982929617,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0129141551218316, 0.00509478070738476,
  0.011615128861512, 0.00472359665186298,
  -0.00419041192306515, 0.00658620539852647,
  -0.0129386930789793, -0.0067787202285608,
  0.00226610473874657, -0.00258396034055602,
  0.0128888664270425, 0.0166854554413789,
  -0.010664068061238, 0.00630742548974073,
  -0.017185155236056, 0.016685455441376,
  0.0172515907719722, -0.00677872022856091,
  -0.00868902553293551, 0.00301709842523676,
  0.00851063250729099, -0.00200794634372106,
  -0.0129386930789792, -0.0067787202285608,
  0.0128888664270423, 0.0166854554413789,
  0.00243775699157289, 0.0040701620543184,
  -4.15781216919734e-18, -0.00677872022856066,
  -0.00414109110299952, -0.00405387918508512,
  0.00614803609105553, -0.00461584648068342,
  0, 0,
  0, 0,
  0, 0,
  -0.000292101678794301, -0.000378144158251909,
  0.000292101678794294, -0.000378144158251909,
  -0.00513459927890502, -0.00202565766784812,
  0.0101699859397645, 0.00542905693934084,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00551537706459859, -0.0055945740186511,
  0.00332734483590391, -0.0107105213165065,
  -3.62832425353654e-19, -0.00694396581485615,
  -0.0128461756510002, -0.00105678586136096,
  0.00774307178261848, 0.000636980919899999,
  0, 0,
  0.00291043790266171, 0.00203943100843179,
  0.017067183458099, 0.0166104692061268,
  0.00526131064823335, 0.00228777342014744,
  0, 0,
  -0.0095214440589286, 0.00287192553461732,
  0.0128610831613167, -0.00694396581485665,
  0.0171121760731734, 0.00379539517610625,
  0.00123121135618336, 0.000541089685905216,
  0.0118777343522401, 0.000937495761427903,
  -0.00914646611402904, -0.00275882202550601,
  0.00525980688457204, -0.00608583458008646,
  -0.00169326675952542, -0.00529994810883636,
  -0.00422448229811054, -0.00413504443621857,
  -0.00858352738557509, -0.0127869471131095,
  0.00858352738557499, -0.0127869471131094,
  -0.00858352738557499, -0.0127869471131095,
  0.00426679586452464, 0.0166104692061374,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000143232926297836, -0.000290811144572189,
  -0.00111194647185847, 0.0035577861601806,
  -0.00385563024391429, 0.0111090542118182,
  -0.00846264749154552, 0.0171820283697373,
  0.0126939712373174, 0.0171820283697457,
  0, 0,
  0, 0,
  0.00424877883130796, 1.38777878078145e-16,
  0.00122489492213495, 0.00365509869602115,
  0, 0,
  0, 0,
  -0.008497557662616, 1.94289029309402e-16,
  0.00726003740413619, 0.011145391268562,
  -0.00247185939786094, -0.00153588005558078,
  0.00423132374577283, 0.0171820283697332,
  1.72786625342116e-17, 0.0109973700354805,
  0.00242237894141986, 0.000947434884715104,
  -0.00562888904922771, 0.00206215032034779,
  0.00424877883130781, 1.38777878078145e-16,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00173426890140546, -0.00169627671044981,
  -0.0126734769710066, -0.0118004889421499,
  0.00421111983988165, 9.43689570931383e-16,
  0, 0,
  -0.00193413465411329, 0.0018009055171489,
  -0.00737714978721344, 0.00785616778334619,
  0.00872298006662178, 0.00286128682242354,
  0, 0,
  0, 0,
  -0.012590822291004, 0.0123149983260296,
  0.00421111983988161, 9.43689570931383e-16,
  0, 0,
  0, 0,
  0, 0,
  -0.00949031040926049, -0.00311298431353368,
  -0.00421111983988182, 9.43689570931383e-16,
  0.0167877630546726, 0.0123149983260592,
  4.12767341006968e-18, 0.0123149983260119,
  0.00328253328372287, 0.0100100772156465,
  0.00119800747253229, 0.000836613778006867,
  -0.00108168334720727, -0.000793490387417217,
  -4.55507421398937e-18, -0.00534503526888891,
  -0.00421727393429834, -0.00534503526888758,
  0.00571041367174591, -0.00219596431331481,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00878706970083128, -0.00162445393560862,
  0.012261138440162, 0.0105484967726059,
  0.00169001144644352, 0.000964928412209187,
  0, 0,
  0, 0,
  -0.000245991584027653, 0.000239989223635273,
  -0.00209007390025115, 0.00605124060639212,
  -0.0041484862597447, 0.0150966301067709,
  0.00416821557364476, -4.9960036108132e-16,
  0, 0,
  0, 0,
  -0.00188348946447243, 0.00153466641679123,
  -0.0122611384401621, 0.0105484967726056,
  0.0124997953501135, 0.00127480779822425,
  -0.0027866747970598, 0.00445899303798464,
  0.0016900114464435, 0.000964928412209187,
  0, 0,
  0, 0,
  -0.00440895265277612, -0.00147650293210533,
  0.0066385793381182, 0.00884384973597374,
  -0.00417158106549998, -0.00257523327570303,
  0.00829697251948943, 0.0150966301067645,
  0.00649671453783371, 0.0101122559250755,
  0.00276971969660288, 0.00282640184770944,
  0, 0,
  -2.86868605206531e-18, -0.00257523327570236,
  0.000498149279305766, -0.000453199970831375,
  -0.00416821557364461, -4.9960036108132e-16,
  0.0165939450389805, 0.0150966301067132,
  -8.26646931815082e-17, 0.0150966301067744,
  -0.00414848625974547, 0.0150966301067508,
  0.0125046467209344, -3.44169137633799e-15,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00285182404479585, -0.000798862115728993,
  -0.0165546649286547, -0.0130224402011854,
  0.00461807737670166, 0.00211395456415736,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000913282948825395, 0.000718418200494619,
  -0.016454220149849, 0.00460920902380357,
  0.00412011952520466, -5.55111512312578e-17,
  0, 0,
  0, 0,
  0, 0,
  -0.00144991279118003, 0.0015207316851123,
  -0.012308390640217, 0.0119925264068098,
  0.00835993486843393, 0.00291409426801104,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.012360358575614, -4.9960036108132e-16,
  0.0123849256038717, -0.00566927919812343,
  -0.0123406651123867, 0.00460920902380485,
  0.0123083906402169, 0.0119925264068093,
  0.00461807737670163, 0.00211395456415736,
  0, 0,
  0, 0,
  -0.00541343208768655, -0.0050358554829214,
  0.00779174671967012, -0.00771328901066998,
  -0.00412011952520449, -5.55111512312578e-17,
  0.00410279688007244, 0.0119925264068107,
  0.0165132341384964, -0.00566927919812449,
  -9.12772654819394e-18, -0.00566927919812271,
  -0.0123654735499271, -0.00106612989962074,
  -0.00413866623216439, -0.0130224402011822,
  0.012360358575614, -4.9960036108132e-16,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00406689166219798, 7.21644966006352e-16,
  0.0121918960393426, 0.00187409655128029,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00338039630242794, 0.00327466449811992,
  0.0121549258921624, 0.00963664043869844,
  -7.54808084264558e-18, 0.00187409655127474,
  0.000355762345904977, 0.000342227976523446,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00230559637677164, 0.00182144852087324,
  -0.00788784007145033, 0.00972105924960304,
  0.0156106458293988, 0.00237277048284901,
  0.000355762345904984, 0.000342227976523446,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00230559637677164, 0.00182144852087324,
  3.16369116573055e-17, 0.00963664043868756,
  -0.0039742441233709, 0.0039044186730105,
  -0.0149777219808815, 0.0101175331045105,
  -0.0121161858454884, 0.0175593708532646,
  0.0122744222318846, -0.0157432838025867,
  0.0121549258921624, 0.00963664043869844,
  0, 0,
  0, 0,
  -0.00161887149785159, -0.000962602488054853,
  -0.0163183057177241, -0.00801580068789226,
  -0.0040795764294307, -0.00801580068791452,
  0.00807745723033043, 0.0175593708528859,
  2.9547100197889e-16, 0.017559370852575,
  0.00260031802926308, 0.00699110228128369,
  -0.00741753971204458, -0.00481790185178149,
  0.00455850831017053, 0.000819558263183362,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00160099793012005, 0.000961084411438218,
  0.0029976386549453, 0.00359898501827094,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00026817099659724, -0.000273228314539742,
  0.000416279714651338, -0.000848260298499881,
  -0.000268170996597236, -0.000273228314539742,
  -0.00272732738486918, -0.00690631563856753,
  0.0159213287515675, 0.0162215820322427,
  0.00577530861868623, 0.00317301989818958,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00326948589309568, 0.00827920464510934,
  -0.0159213287515662, 0.0162215820322454,
  -0.00604004306164168, 0.0020664612072479,
  0.00957740026524218, 0.00797899461960194,
  0.0159213287515668, 0.0162215820322427,
  0.00577530861868608, 0.00317301989818958,
  0, 0,
  0, 0,
  -0.00400859835333591, -7.7715611723761e-16,
  0.00805045646140464, -0.00966543187154212,
  -9.34551857129146e-18, -0.00966543187153701,
  -0.0120756846921071, -0.00966543187154817,
  0.0120334524919248, -0.00146483328574293,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00394531228663468, -3.33066907387547e-16,
  0.0118956763527266, -0.0107163746395927,
  0.000193034817869313, -0.00220880385961447,
  -3.72647871779848e-18, 0.0154183802296693,
  1.82849127309958e-17, 0.0069217443594356,
  1.61182257888486e-17, 0.00692174435943549,
  0.00181452137949918, 0.00490390549919256,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00928146180986582, 0.00379699806960943,
  0.00396522545090884, -0.0107163746395922,
  0.0156652739529127, 0.0154183802296343,
  -0.00475193173518506, -0.00105593640120311,
  0.0133600346314453, 0.00314634843526373,
  0, 0,
  0, 0,
  0, 0,
  -0.00333634907773442, 0.000478783560369567,
  -0.0156652739529127, 0.0154183802296315,
  0.00391631848822811, 0.015418380229667,
  0.000635009240959618, -0.000833334840352862,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00120565548236705, 0.000874002030578802,
  -1.51609146990572e-17, 0.00632572644793222,
  0.00195997383915992, 0.00189442853878835,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00195997383915992, 0.00189442853878835,
  -0.00863092839325072, 0.00798881120314043,
  0.00896582457565813, 0.00355436385926744,
  -0.00818244105285707, 0.00567503953733284,
  0.00195997383915991, 0.00189442853878835,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0155084495198686, 7.99360577730113e-15,
  0.0154579749086374, 0.00632572644794432,
  0.000479984551873737, -0.000117398815371705,
  0.0101989521046586, -0.00664174853414606,
  0.00077349877213617, -0.00150738461137528,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00380408368408664, -6.66133814775094e-16,
  0.0113169391661176, 0.0147644927820448,
  0.00181702197624836, 0.00183659817284454,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00143897781394615, 0.00436344313674286,
  -2.12314043277957e-17, 0.00601991889320075,
  -2.89428199162786e-17, 0.00601991889320075,
  -0.00619956324208583, 0.00841157783187318,
  -4.72620482273567e-17, 0.0147644927820664,
  0.00765893040606255, 0.0058762078748068,
  -0.00760816736817295, -1.4432899320127e-15,
  0.0114864309031668, -0.0116101831926377,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00417720739695963, -0.00637973709432604,
  6.5925591562858e-17, -0.0118076721700912,
  0, 0,
  -0.000605974456871958, -0.00239120993337072,
  -2.69543089576658e-17, -0.011807672170091,
  3.83009899053706e-19, -0.0118076721700912,
  -0.00202639107285907, -0.00390829002095872,
  0.00417720739695956, -0.00637973709432615,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00444309389570144, -0.00140787649007468,
  -0.00805050783242756, 0.00764235701032889,
  0.0052050193218004, 0.00233443227090879,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00550464169071157, 0.00153185589437554,
  0.00084004217652136, -0.00110495152293888,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00501441234499813, -0.00388468111955498,
  3.40309084982387e-17, -0.0119987023993136,
  -4.0512986307427e-19, -0.0119987023993136,
  -0.0146904476334602, -0.0119987023993703,
  0.000875877677934657, -0.00116336249994997,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0109556943824648, -0.00331004534215007,
  0.00360920398929466, 0.0143815033134491,
  0.00305540624468121, -0.0011538043989413,
  -0.00446010068816952, 0.00698089000003521,
  -0.00360920398929497, 0.0143815033134795,
  0.00502774571255759, 0.0102102519832529,
  0.00100170660460436, 0.000818162913748255,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00560525995459279, 0.00818099136012074,
  -0.0144368159571795, 0.0143815033133877,
  0.00979772169568103, -0.00713184617720741,
  0.000912797112125942, -0.00181859971499776,
  0, 0,
  0, 0,
  0.000662617609092323, -0.00267052181993233,
  0, 0,
  0, 0,
  0, 0,
  -0.0106708953636815, 8.99280649946377e-15,
  0.0105627840741667, 0.014190258434821,
  2.05445773308734e-16, 0.0141902584347746,
  -0.0070418560494446, 0.0141902584347954,
  0.00711393024245435, 3.99680288865056e-15,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0105627840741675, 0.0141902584348204,
  0.00628532797463536, 0.00139568398186707,
  -0.007086571740064, 0.00543066698977424,
  0.00717533802894369, -0.0121894551917778,
  0.00199544236314448, -0.00426434917410956,
  -5.59817545905376e-05, -0.000433438647556406,
  -1.53189180448044e-17, 0.00543066698976835,
  -0.0105627840741668, 0.0141902584348204,
  0.00748117546417868, 0.00737975800847535,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00802585365013644, 0.00315230460752958,
  0.0106708953636815, 9.10382880192628e-15,
  -4.07822718195711e-17, -0.0121894551917909,
  4.6252792779326e-17, -0.0121894551917909,
  0.0139932226902571, -0.0123798999177256,
  -9.2563117732815e-17, -0.0123798999177278,
  3.63010215013901e-17, -0.0123798999177278,
  5.53472653983936e-17, -0.0123798999177278,
  -0.0104949170176928, -0.012379899917727,
  0.00346166474568418, 0.00153075222676269,
  -0.010284943093596, 0.0139992104755605,
  0.00993787638603214, 0.00850303858919021,
  -0.00993787638603217, 0.00850303858919021,
  0.00993787638603214, 0.00850303858919021,
  0.00151865083909225, 0.00268712158937157,
  0, 0,
  -0.00141618723996789, 0.00167054739604033,
  0.00141618723996789, 0.00167054739604033,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0104949170176932, -0.012379899917727,
  0.00141618723996789, 0.00167054739604033,
  -0.00749779413831142, -0.00226446880763931,
  0.00699661134512864, -0.0123798999177278,
  0.00503316046485311, -0.00381759959161909,
  -0.0103967719010255, 5.55111512312578e-16,
  0.0137132574581276, 0.0139992104755625,
  0.00261314011929375, 0.000694670219275051,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00482706506465837, 0.00171095218464723,
  0.00690350677537808, 0.0052362377139501,
  0.00151865083909224, 0.00268712158937157,
  2.11044427695784e-17, 0.00523623771394988,
  -0.00444617501490231, 0.00999557699189602,
  -0.00999443152483965, 0.0138083865450023,
  -0.00333147717494677, 0.013808386545002,
  0.00999443152483925, 0.013808386545002,
  -0.00768856848593776, 0.00248727796733805,
  0.00999443152483991, 0.013808386545002,
  0.00132082957901941, 0.00162551383173926,
  -0.00673980141445856, -9.99200722162641e-16,
  0.00673980141445856, -9.99200722162641e-16,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.00417776810046657, 0.00987945039566474,
  -0.00417776810046631, 0.00987945039566474,
  0, 0,
  -0.0103816979438754, 0.0042152678820625,
  0.0102138959342067, -0.0125700009908467,
  -0.00490502697080549, -0.00193752762979305,
  0.007526441760178, 0.00296478788070909,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0100679105225821, 0.00504176236068565,
  0.00673980141445857, -9.99200722162641e-16,
  0, 0,
  0, 0,
  0, 0,
  -0.00323968080184071, 0.002762263129089,
  -0.012922143335294, 0.0136178181173302,
  -0.00328184271290032, -0.00407992235581345,
  0.00921608885012094, 0.00825755115799531,
  0.000267620804384906, 0.0011472109520948,
  -0.00637982436570169, -0.00636709767662214,
  0.00981004427284759, 0,
  0, 0,
  -0.00122761943443942, 0.00157899379365556,
  0.00122761943443944, 0.00157899379365556,
  -0.00449199018246877, -0.00668716143989945,
  0.00345309734895174, -0.00918945260404613,
  1.53560656686399e-17, -0.00407992235581345,
  -0.0040972924333685, -0.00711129354355378,
  4.23965485847334e-17, -0.0127597168359771,
  0.00398746809512247, -0.00197869554513574,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00122761943443939, 0.00157899379365556,
  -0.00969160750147042, 0.01361781811733,
  -2.5627461877473e-17, 0.0136178181173303,
  -0.012922143335294, 0.0136178181173302,
  0.00654002951523183, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00130858718097232, 0.00252470469990074,
  -0.00651210895015769, 0.00484724165625683,
  0.00654002951523175, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000859452008728341, 0.0034725949342983,
  -0.00427604055761685, 0.00754661349195274,
  7.64679853092567e-17, 0.0134275419936013,
  0.00113675367582437, 0.00153100852485966,
  -0.00415492005328365, 0.00186100014944135,
  -1.06118528036353e-16, 0.0134275419936005,
  0.00305469987846585, 0.00271671536669504,
  0, 0,
  0, 0,
  0, 0,
  -0.00700109879121594, 0.00277002082142697,
  0.00312561478508461, 0.0134275419935996,
  0.00113675367582437, 0.00153100852485966,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00120817733810893, 0.00244080557229642,
  -2.46813970457283e-17, 0.00465267628547472,
  -0.00937684435525412, 0.0134275419935894,
  0.00407253409399188, -0.00437525654974058,
  -0.00215158325096603, 0.00024476996280054,
  0.00633211492499135, -1.33226762955019e-15,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00113675367582438, 0.00153100852485966,
  -0.00312561478508451, 0.0134275419935986,
  0.0093768443552544, 0.0134275419935912,
  -0.00937684435525346, 0.0134275419935894,
  0.00640964066255223, -0.0129489985883,
  -4.87028994363108e-17, -0.0129489985882952,
  8.89616499994726e-17, -0.0129489985882953,
  0.00285176847577018, -0.0026189932509606,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00104842005945796, 0.0014815788413588,
  -5.53851356106272e-17, 0.0132376015234658,
  0.00186789842211345, 0.0051415420552301,
  -1.21959474523771e-17, 0.00445806690411721,
  0.000661639402129612, 0.000701248700338164,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00287295518014068, 0.00266852502826032,
  -0.0120673735492774, 0.0132376015234951,
  0.0122326344543857, 7.21644966006352e-15,
  -0.0122326344543862, 7.21644966006352e-15,
  0.00611631722719306, 1.22124532708767e-15,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000661639402129624, 0.000701248700338164,
  0.00111106897049472, 0.00235516708659655,
  -0.00194427448958461, 0.00166712641560496,
  -0.00611667027365806, -1.81852197641552e-05,
  0.00671963736217403, 0.00266551740434018,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00383049295777613, 0.00438025323677504,
  0.0117858118583641, -1.86517468137026e-14,
  -0.0117858118583647, -1.86517468137026e-14,
  0.00371482339402064, 0.00194576050868023,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00653164462050131, -0.00259985962975928,
  0.00580871151380499, 0.013048048172817,
  -7.57827587056103e-17, 0.0130480481728299,
  -0.00293277092632075, 0.00426341415334441,
  0.00322446877089961, 0.00936934207141815,
  0.000609163774493332, 0.000678917180563454,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.00394977710582304, 0.00671943946821663,
  -0.00617042882718024, 0.00246508097220299,
  0.0111531624240472, 0.0128589435587592,
  0.00167584039712894, 0.00478710385601511,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00439902734957566, 0.00374185646462499,
  -0.00557658121202392, 0.0128589435587738,
  0.00865131318130871, -0.00427554930916685,
  -0.00102801338006398, -0.0015803190197623,
  -0.00578306889948857, -0.00693841435110021,
  0, 0,
  0, 0,
  -0.00199414087216559, -0.000715573131124358,
  0.00385707999252066, -0.00777218047324468,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00837346310132109, -0.00419196359878327,
  0.00736817053719761, 0.00758399322173853,
  -0.00736817053719761, 0.00758399322173908,
  0.00788353610690289, 0.004592960196528,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000785719440281405, -0.00373028444385437,
  0.00102734823633816, -0.001625814062019,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000800348970158289, 0.00132482536795087,
  0.00059068487811491, 0.00293329912389417,
  -0.00542436831169435, 2.22044604925031e-16,
  -0.00334636278073254, 0.00698446396985963,
  -0.0106751643041182, 0.0126703621221984,
  0.00366890413169696, -0.00175538866817837,
  0, 0,
  -0.00263855264101404, -0.0138864203340634,
  0.00333479537152771, -0.00992716234868896,
  0.000638448480644053, -0.000782536491255259,
  9.45868718288956e-17, -0.00522223565232283,
  -4.89232805474002e-17, -0.00522223565232283,
  1.04523009797279e-17, -0.00522223565232283,
  0.000638448480644037, -0.000782536491255259,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000638448480644022, -0.000782536491255259,
  -3.14859436920198e-17, -0.00522223565232283,
  -0.0037860684570688, -0.00789304039045169,
  -0.0105542105640548, -0.0138864203340917,
  0.00517982781058955, -8.88178419700125e-16,
  -0.000723832783571169, 0.00126981817329186,
  -0.00763801370083095, 0.0124823946860918,
  0.00259549135931595, -0.00156036281572536,
  -0.00254600456694379, 0.0124823946860989,
  0.00773108126729843, 0.00367920226153817,
  0.000723832783571175, 0.00126981817329186,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0103596556211797, -5.99520433297585e-15,
  0.00517982781058971, -8.88178419700125e-16,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00582452585139522, -0.00305539690946,
  0.00102172596318104, -0.00166975174868833,
  -0.00559227519755634, 0.00225375742448841,
  0.00517982781058956, -8.88178419700125e-16,
  -0.00102172596318104, -0.00166975174868833,
  0.00248393357130878, -0.00541033943195435,
  -1.5332080240294e-16, 0.0122951532618956,
  2.56577669327368e-17, 0.0122951532618955,
  -0.0072602476907122, 0.0122951532619094,
  0.00251496557688618, -0.0140713780671331,
  0.00347122665673471, -0.00164430976101648,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00160248817691755, 0.000872608377390782,
  -0.0096803302542834, 0.0122951532619318,
  0.00492884471823117, 1.88737914186277e-15,
  0, 0,
  -0.00202064681493636, 0.00239028347269665,
  -0.00968033025428353, 0.0122951532619318,
  0.00225325596727607, -0.00940847700399039,
  7.86580383414557e-17, -0.00194426700859307,
  -0.00242008256357067, 0.012295153261898,
  0.00490381349247493, 0.0034843828375124,
  0.000679963417974113, 0.00190221735320795,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000630121326931674, -0.000800327890133956,
  4.54764607138499e-17, -0.00541033943195546,
  -2.49399329622714e-16, -0.0140713780671368,
  -0.0100598623075443, -0.0140713780670814,
  0.00502993115377115, -0.0140713780671272,
  0.00187235986768468, -0.000665198482630691,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00101099034186899, -0.0017121015327709,
  1.29927099110329e-16, -0.0140713780671368,
  -0.0100598623075418, -0.0140713780670814,
  0.00502993115377173, -0.0140713780671272,
  0.00400124378286146, -0.00127034380164925,
  0.000650644624201813, 0.00121346478571416,
  -0.00777121809001213, -0.00399845176035474,
  0.00458236091943618, 0.0121087776460511,
  1.04667589522243e-16, 0.0121087776460491,
  0, 0,
  0, 0,
  -0.00477406245340082, 0.00290849015907924,
  0.00693369212673233, -0.00866354292511762,
  -9.03558433648573e-17, -0.0055974880922951,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000421446273158443, 0.00251552228732677,
  -0.0068735413791538, 0.0121087776460529,
  0.00693369212673228, -0.00866354292511762,
  0.00107262824232154, -0.00283439412815656,
  0, 0,
  -0.00934346694820214, 2.66453525910038e-15,
  -0.00229118045971811, 0.012108777646052,
  0.00368717876043425, -0.00513174792446969,
  1.01810380420159e-17, 0.00328952379507053,
  1.00568790415035e-17, 0.00328952379507053,
  -0.00929508753075096, 0.00328952379507275,
  0.009164721838872, 0.0121087776460584,
  0.00271337134590523, 0.00653973522903883,
  0.000580914090293459, 0.00115578381257153,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00180353933100556, -0.000638271078681196,
  -9.45215752265516e-17, -0.0142551286090827,
  -0.00238827970475924, -0.014255128609083,
  0.00916472183887213, 0.0121087776460584,
  0.00149351841541906, 0.000886894480210509,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000618558371245166, -0.000817262750598902,
  -0.00693369212673218, -0.00866354292511751,
  0.00311028592883823, -0.00422213034215568,
  -0.000618558371245156, -0.000817262750598902,
  -0.00942609491035261, -0.00559748809229088,
  0.000514760668141599, 0.00109679357719683,
  0, 0,
  0, 0,
  0, 0,
  -0.000330615554481339, 0.000528328559929125,
  -0.00438556299405258, 0.00309462624885093,
  0.0043189147638336, 0.0119234446382628,
  -8.05133724686209e-17, 0.0119234446382668,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000535085557106855, 0.00171014931386759,
  -5.25025703643511e-17, 0.00309462624885204,
  3.16747159200171e-17, 0.00309462624885204,
  -5.28344646698646e-17, 0.00309462624885204,
  4.22545902949408e-17, 0.00309462624885204,
  -4.22545902949408e-17, 0.00309462624885204,
  0.00677595334863899, -0.0144374319409739,
  0.00323122262140398, -0.00152005209724848,
  -0.00259975560201812, 0.00675393163898219,
  -9.38341788717892e-17, 0.0119234446382663,
  2.61832105589011e-17, 0.0119234446382668,
  -0.00647837214575071, 0.0119234446382586,
  0.00215945738191689, 0.0119234446382654,
  3.27290131986264e-19, 0.0119234446382663,
  0.000907046286064018, 0.00226274661566395,
  0.00037138763076317, 0.00237393177032308,
  0, 0,
  0, 0,
  -0.000371387630763154, 0.00237393177032308,
  -0.00215945738191706, 0.011923444638265,
  0.00647837214575084, 0.0119234446382595,
  3.27290131986264e-19, 0.0119234446382663,
  0, 0.0119234446382668,
  0.00037138763076316, 0.00237393177032308,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00225865111621275, -0.0144374319409601,
  0.00881763321511236, -6.66133814775094e-15,
  0, 0,
  0, 0,
  0, 0,
  -0.00428314292918507, -0.00302235461085032,
  0.00351885546213789, -0.00822585999648862,
  -0.00482246167657597, -0.00758082318310582,
  0.00647837214575102, 0.0119234446382595,
  -0.00215945738191668, 0.011923444638265,
  -0.00225865111621275, -0.0144374319409601,
  -0.00215945738191631, 0.0119234446382595,
  0.000946662134789845, -0.00182926921718707,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00675008364160819, -0.00363576218194628,
  0.00414042449626523, 3.5527136788005e-15,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00112734482782646, 0.00371040978396708,
  2.76957836443694e-17, 0.0117393811821811,
  0.000452293658948756, 0.00103651215953104,
  0, 0,
  0, 0,
  0, 0,
  -0.000468918378005127, 0.00161191603401978,
  -0.00189812549482838, 0.00835975967418601,
  -2.83712905625248e-17, 0.0117393811821811,
  2.76957836443694e-17, 0.0117393811821811,
  0.00460004254146114, -0.00769634492276805,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00029120492114197, 0.000500511286816163,
  0.000468918378005148, 0.00161191603401978,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -5.01354682898718e-17, 0.0117393811821811,
  -0.00810030406066505, 0.0117393811822448,
  0.00837263547397522, -0.00596813481221226,
  -2.11403901246517e-17, -0.00596813481224445,
  -0.00147048574638969, -0.00647634072542025,
  -1.31584566792191e-16, -0.0146179793769818,
  0.00173506037191855, 0.00169301227826701,
  -0.00405015203033233, 0.0117393811821918,
  0.00195574315463275, 0.00477496112932374,
  0.000468918378005105, 0.00161191603401978,
  -0.000291204921141939, 0.000500511286816163,
  -0.00823639364562078, 0.00289969158663372,
  0.00810030406066505, 0.0117393811822439,
  -0.00810030406066505, 0.0117393811822448,
  -0.00212623952939095, -0.0146179793769334,
  0.00398241618434546, -0.0147963671545421,
  0.00140295134541891, -0.00663428691530799,
  0.000914075427099459, -0.00186488889317316,
  0, 0,
  0, 0,
  -0.00208229086154906, 0.00372228567060229,
  -0.00180336175571491, 0.00100892829493548,
  0.00225868359234466, -0.00298153518956212,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.000726638402465082, -0.00444744442067768,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00294772336154939, -0.00138208189886524,
  0.00377640486902417, 0.0115568835255062,
  0.00104025423415157, 0.00352927580991103,
  0.00566460730353651, 0.0115568835254858,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00208229086154911, 0.00372228567060229,
  -7.356908119047e-17, 0.0115568835255224,
  0.00212914369042918, 0.0060800395785312,
  -0.0010402542341515, 0.00352927580991103,
  -0.00755280973804885, 0.0115568835254249,
  0.00755280973804777, 0.0115568835254249,
  6.96067456180318e-17, 0.0115568835255224,
  -2.87755338193558e-17, 0.0115568835255224,
  0.0021291436904293, 0.0060800395785312,
  0.000393612123491167, 0.000974957450621705,
  -0.000393612123491137, 0.000974957450621705,
  -0.00576866756170231, 0.00270472159007928,
  0.00353889456351453, 0.00528257803391141,
  0, 0,
  0, 0,
  0, 0,
  -0.00208229086154911, 0.00372228567060229,
  0.0018882024345122, 0.0115568835255162,
  -0.00104025423415159, 0.00352927580991103,
  7.356908119047e-17, 0.0115568835255224,
  -0.00566460730353649, 0.0115568835254858,
  0.0079648323686879, -0.0147963671543905,
  -0.00796483236869115, -0.014796367154531,
  0.00554125970967245, -0.00964295227515333,
  0.000644414872197302, -0.00103389813021981,
  0, 0,
  0, 0,
  -0.0018884153377872, 0.00394253425997082,
  0.00187338290898736, 0.00394927352602936,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.000844724704651204, 0.0102765415842283,
  0.000168885631940187, 0.00186231228092626,
  0.00271522007239858, -0.008222423340976,
  0.000566187572591348, -0.0027144322683077,
  -4.52354051567755e-05, -0.00019034517921579,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000338804844956307, 0.000912147229081173,
  0.00150986266037736, 0.00800736514281142,
  -4.8008547072416e-17, 0.0025097186127816,
  0.0003388048449563, 0.000912147229087168,
  -0.000940683208056534, -0.00187445940239717,
  0.00700742833714565, -0.00448003401934693,
  0.000588525835263779, -0.0057225832664427,
  0.00103732783319822, -0.00219117424809157,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00168073982978148, -0.000711558969864967,
  -0.00744475129987076, -0.0142069425665385,
  0.00735556236162567, -0.0115966870461444,
  0.000110433465064725, -0.011437331956218,
  0.001816679851382, -0.00317660128959663,
  0, 0,
  0, 0,
  0, 0,
  -0.00159662500889728, 0.00188427300828531,
  -0.0075434613793661, 0.0129188041085677,
  0.00319379239740904, 0.00919850673442757,
  0.000828741218468624, 0.000979773442979504,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00163255326719347, 0.00582083131283428,
  -4.31774103056794e-05, 0.0104820071337728,
  -0.00543335768588079, 0.0104171006149736,
  0.0036085515880336, -0.00404313567523928,
  0.000364920565111779, -0.00609184802203266,
  9.4387838174449e-06, -0.00643076386379904,
  6.67275772831764e-06, -0.00638283191897182,
  -0.00546193674013951, -0.00637160366133149,
  0.00476705582186331, -0.00992244012455545,
  0.000430322541228437, -0.000664651981238773,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000783511317614848, -0.00284985087290823,
  -0.00746582898437026, -0.00761803427293239,
  0.00650140843054674, -0.00857003221700769,
  -0.0047870539893637, -0.00545135889911674,
  0.000133063009186382, -0.00851807714615838,
  -8.93538019011241e-06, -0.000985698382722777,
  -0.000495700885878455, -0.00194971287128709,
  0.000323856731081269, -0.000739658414153022,
  -9.36519455295419e-05, -0.000222822000980338,
  6.12037576932765e-06, -1.38478925080232e-05,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000424256033762618, -0.000609517927039338,
  -4.13495382506999e-05, -0.00720340733555025,
  -0.00146254054685843, -0.0137330583756277,
  -0.00337242456186277, -0.0159864045394733,
  0.00533569355967917, 0.00891926061662374,
  0.00135352711743652, 0.00247923787948956,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -5.52159715678961e-05, -0.000136389593399899,
  -0.000526862570113897, -0.00339419107703831,
  0.000829598185649071, -0.00326614445901718,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  3.38183527755659e-05, -0.000152721381964538,
  -3.26976401338611e-05, 5.11940944376565e-05,
  -0.00429069311599927, -0.000845773787852444,
  0.00243257214024085, 0.00735381141364799,
  -0.000301925139246219, 0.0100607146046932,
  0.00167776323494203, 0.0009665593898045,
  0, 0,
  1.9136447831977e-05, -0.00139645876336902,
  -0.00116514890932819, -0.00727636423595701,
  -0.00798142781565031, -0.0136721088504996,
  0.00424887195676673, -0.00684804744168654,
  4.38883139945187e-06, -2.6719577850276e-06,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00100943726795703, 0.00158468559853198,
  -0.00402975165325958, 0.00898365481073249,
  0.00136458727461585, -0.0110887780928439,
  0.00135936982734438, -0.00671197515212452,
  0.000224142801648697, -0.00383448239816486,
  0, 0,
  -5.98835343766687e-06, -1.49756732019668e-05,
  -0.00013137588163006, -0.000917756798652469,
  -0.000963025115007651, -0.00718775506118674,
  -0.000351798546044883, -0.0108553690937592,
  -0.000494550935200934, -0.0123495163815637,
  -0.00643238432615786, -0.0124344843103175,
  0.00777778462429294, -0.0117769544223778,
  -0.00341954605015741, -0.00736314088470769,
  -0.00546339010262912, -0.0173721399885658,
  -0.00260176688923595, -0.0101331084275997,
  0.00239040843960591, -0.0149728154434321,
  0.00216443879063491, -0.000217969327680034,
  0.000888803161862256, -0.00604942667410113,
  -0.000780643605729729, -0.00695408304219658,
  -0.000863682873843487, -0.00973241300937144,
  0.00100184398578411, 0.000732826394797659,
  -4.72614403235654e-05, -0.000114276454790119,
  6.92228384337606e-05, -0.00422091059544005,
  0.000347058173541218, -0.00131479983713811,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  4.27104211997497e-05, -0.000679843018314585,
  5.98835343769223e-06, -1.49756731999684e-05,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -4.79235840811066e-06, -1.25581031795718e-05,
  1.54610067711035e-05, -3.99250444713672e-05,
  0, 0,
  -0.000352076983671567, -0.000653979463911103,
  3.73352473793496e-05, -0.00712879282134926,
  2.68277308875959e-05, -0.00691323976129055,
  1.56831074226438e-05, -0.00676971857324249,
  -0.00267807524186808, -0.0108115357556517,
  0.00220939806594992, -0.00775176427307467,
  -1.56831074224785e-05, -0.00676971857325759,
  -2.68277308876583e-05, -0.00691323976131142,
  -0.0033014863734771, -0.00939649655917618,
  -0.00126127745210768, -0.015902742139009,
  0.00286831546120353, -0.0105740077842771,
  -0.000177006099776004, -0.0106455750545749,
  0.000328291779810733, -0.00438952387952085,
  4.97957297589554e-05, -0.000126657208286529,
  0, 0,
  -5.98835343766676e-06, -1.49756731999684e-05,
  -0.000131375881630136, -0.000917756798638925,
  -0.000153934557192198, -0.00241537202827224,
  -0.000187175647631084, -0.00401294403275343,
  -0.000227677457179058, -0.00570929598088177,
  -0.000290736807945472, -0.00750628940105247,
  -0.00038376058938833, -0.00940177817374432,
  8.28973378979535e-05, -0.011060336328544,
  -0.000378559596687847, -0.00769418220765861,
  0.000542085830883195, -0.00629957639878431,
  0.000381165104066049, -0.00593062323955507,
  -0.000415554940317957, -0.005023105790956,
  0.000424996070039736, -0.00608225288630271,
  -0.000627015170090644, -0.00730568602880788,
  -0.000468513205603576, -0.00955295128927292,
  0.000278088299688812, 0.00619406276611167,
  0.000732906726236582, 0.00452155835139822,
  -0.000971295233614356, 0.00556315273721841,
  0.000217604137674572, 0.00100110705367262,
  7.75575966474358e-05, -0.0046386436496193,
  0.000250035993968764, -0.00527209555292818,
  0.00041931561699302, -0.00241863881642979,
  -6.01998290279258e-05, -0.00102376929503323,
  0.00015822574202351, -0.000779972795028394,
  0, 0,
  -0.0010296609177796, -0.00331817624777697,
  -0.0013238644327347, -0.00881002214908078,
  0.00219928677656259, 0.00734111123249037,
  0.000222697795729636, 0.000278901573459889,
  -0.00206171824940451, 0.00577074408050327,
  -0.000286350506870248, 0.0110655830487529,
  0.00153703860110465, 0.0036751150921126,
  0, 0,
  -1.42133966238287e-05, -4.47812819057702e-05,
  -0.000710661048228714, -0.00223773048490039,
  -0.00748963442360429, -0.00483957116173639,
  0.00194102030013486, 0.00631919176152884,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -7.30332326535471e-06, 1.84733164168005e-05,
  -0.00122980159544064, 0.00520061756861523,
  -9.2892995463933e-05, 0.00945134154403204,
  -0.00272368907406685, 0.00938721746511351,
  0.00679013437826879, -0.0162591153820297,
  -0.00104841083096333, -0.0154678149230902,
  -0.00365161036343202, -0.0166857664614855,
  0.00565422889473945, -0.000678780904341814,
  0.00022659760773274, 0.000828944717992774,
  -0.00628433990547639, 0.00563415386597765,
  0.00431833855634853, -0.00905378793163836,
  0.000944802284987324, -0.00248678552729942,
  -7.40047832192739e-05, -1.80650364918211e-05,
  -0.00534333418801613, 0.000320722896069769,
  0.00357401590180454, -0.00220247463511369,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000631805335775029, -0.000824965330605387,
  -0.00697016439577183, -0.0127115568124836,
  0.00228441499850375, -0.00780732973918496,
  0.000211331336088578, -0.00775110591513695,
  0.00016380235315925, -0.00639078341950827,
  0.000137321869372455, -0.00514464234271395,
  0.000109032158088041, -0.00400659604978926,
  9.42225101927933e-05, -0.00297897954473569,
  -0.000197031287173029, -0.00283686694659901,
  -0.000685468607204447, -0.0101531151495435,
  0.00508345657082608, -0.0171969769496541,
  0.00124052717470387, -0.0167512104910041,
  -0.00058971480021851, -0.0163729361693823,
  0.00538831948556556, -0.00773922317473819,
  -0.00275016855365135, -0.00598903683225527,
  0.000284332340138321, -0.0145180654004573,
  -0.00104841083096127, -0.0154678149279313,
  -0.00365161036343895, -0.0166857664621543,
  0.00662356491834756, 0.00727610934690204,
  0.000932873418839189, 0.00853189460692194,
  -0.000550529321419588, 0.00652356878718252,
  0.00156059866570837, 0.00634462170397732,
  3.17146152943035e-05, 7.53136883278049e-05,
  0, 0,
  0, 0,
  0, 0,
  -0.000105241197128862, -0.000288595683189952,
  -0.00491323498724057, -0.00827842172278404,
  0.00160688407454704, 0.0167213779472943,
  0.000113187621264233, 0.0109192229047748,
  0.000982009946526235, 0.00231925158800683,
  -0.00134714644910181, -0.00101053551027586,
  -0.00474772416468565, -0.0122090378422046,
  0.00212563517364749, 0.00143345965287289,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -9.03672242953927e-05, -0.000270090172909132,
  -0.00103175151688617, -0.00647895604942161,
  -0.00343595483515873, -0.0118316477321847,
  -0.00351611446682037, -0.0174678918285847,
  0.00669257297534226, 0.0139768301174312,
  0.000600119464859158, 0.000926029871530565,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -8.02025872040854e-05, 0.000285534890753558,
  -0.00440875799214343, -0.00123175543005449,
  0.0063640125320379, -0.0184623444480683,
  0.0022826443426396, -0.00430446159199249,
  -0.00136993043315131, 0.00312903528980213,
  -0.00488976715568001, 0.014783723210275,
  0.00386565583408914, -0.0143834328918686,
  0.000177057409019423, -0.012580425836157,
  -0.00618266141327548, -0.0168402833801575,
  0.0041510996655302, -0.0163467134483646,
  0.000454383675857927, -0.0158716237217018,
  -4.93281814073718e-05, -0.00522975051919894,
  -0.00012846410136525, -0.00582016457008594,
  0.000479753926609761, -0.00480810431112633,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00088879306916513, -0.00406076629949514,
  6.57044158548037e-05, -0.00634861018641608,
  -0.000746514939645457, -0.0110625378706259,
  0.00103704424977933, -0.0145161512400316,
  0.000602216611436202, -0.0118968362431395,
  0.000356233609404819, -0.00951066976977244,
  -0.00254598669720107, -0.0155459307081303,
  0.00527181561679038, 0.0193872133572719,
  -0.000285371026265356, 0.0114509577240762,
  -0.000315113638368711, 0.0128164084875726,
  -0.000389472946446404, 0.0140569007730413,
  -0.000475599831956984, 0.0151579003064948,
  -0.00423381925115061, 0.0154975051043789,
  0.00617904932961334, -0.00490519216493057,
  0.000840140945895105, -0.00546110181891302,
  7.43844406154957e-05, -0.00356346276300346,
  0.000191727842321888, -0.00669902603512185,
  -0.000878112013382769, -0.00728792494523067,
  0.000308774822148763, -0.0145575004921079,
  0.000801645891109533, -0.014539811164735,
  0.000811189327332954, -0.0118516726418025,
  -2.92828252936895e-05, -0.00740427606538274,
  -0.00415923934341517, -0.000840257495211105,
  0.00211367018828609, -0.0157956433173563,
  -4.93281814075232e-05, -0.00522975051919539,
  9.2840774554641e-05, -0.00522574941103571,
  8.75627937189769e-06, -0.00367091903020289,
  -0.00360291129550956, 0.00334047403049054,
  0.00475297030466791, -0.00798172878788161,
  -0.000166500928201467, -0.00984397128381542,
  0.000408049288952371, -0.00846639610329603,
  -7.79688496485145e-05, -0.0090570663288212,
  -0.00020161038689874, -0.0109942930247866,
  -0.004235377830955, -0.015660242199135,
  0.00362942288494244, 0.00800828711775559,
  1.66628364280746e-05, 4.60811223972346e-05,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00256177750186104, -0.00170359088970629,
  0.0056965117880686, -0.0174982355751676,
  0.00255266413587011, -0.0153466008571901,
  0.00084207728290073, -0.00320305718034986,
  -0.000684575798704722, 0.00284773584996856,
  -0.000642529893503288, 0.00876258978729338,
  -0.00121384696822152, 0.0117450067256717,
  -0.00512683211908724, 0.00706357101955635,
  0.00555329687528192, -0.0172616529238867,
  0.000738867290358484, -0.00890890401414501,
  0.000445932746085554, -0.00726018154452035,
  -0.000370212228663027, -0.00373851665064517,
  0.00024649572104425, -0.00256593189680876,
  -0.000140997757293974, -0.00306515877687508,
  5.67690786475257e-05, -0.00022290068988795,
  0, 0,
  0, 0,
  0, 0,
  -0.000331263596770703, 0.000318713187604125,
  -0.00231700182500134, 0.00126463517236242,
  -0.0053063265251342, 0.00125331502413495,
  0.00551841960553538, 0.000579924875818927,
  0.000343162691411488, -0.00826075656450076,
  0.000171525643534853, -0.00701279909194974,
  7.3796024098262e-05, -0.0057597804293692,
  -0.000492306673691799, -0.0126725913084349,
  0.000219306649618938, -0.0115773722656429,
  -0.00496005909641118, -0.01713082102762,
  0.00502574851288146, 0.010778027337937,
  0.00098538680316057, 0.00829645512864197,
  0.000117103253027605, 0.0106224892235001,
  -0.000254417207665492, 0.00276666797125724,
  0.000911253308977942, 0.000148068248302158,
  -5.93137372061917e-05, -0.00142592687905241,
  -0.000222940692443254, -0.000377801404271239,
  -0.000477207429606843, 0.0025801979682345,
  -2.10000751462629e-05, 0.00934586329853948,
  -8.71876781304908e-05, 0.0103089753267653,
  4.89463038420551e-05, 0.00249447725900653,
  -0.00111541036036166, 0.0118781269321582,
  0.000366425200736654, 0.0141502268243419,
  0.00130697147180954, 0.00230690390291199,
  7.78763112629677e-05, 0.000254516519540449,
  5.38834861238395e-05, 0.00234409844836669,
  1.52386870830509e-05, 0.00185469345475231,
  -0.000801743394107532, 0.000821945010448299,
  -0.00468810046218524, 0.000819856911883354,
  0.00409555570625849, 0.0202988793695511,
  -0.000266399986170179, 0.0164218407466052,
  0.000353150517263142, 0.0131278798713073,
  0.00178578877080807, 0.014296292309635,
  0.000731724658264168, 0.00826308727016789,
  0.000155074710959364, 0.000524009619452759,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00107132992005573, 0.00317445219310963,
  -0.00192649071700691, 0.00820329400281783,
  0.00324690143205257, 0.0113938645543228,
  0.00125946489489472, 0.00213055619453595,
  0.000115477762796425, 0.00298380243729301,
  -0.00103845863751038, 0.0101463038068068,
  0.000215061323906496, 0.00881608307564474,
  -0.00399740661680044, 0.0197264785191935,
  0.0049465918660459, -0.0176618264750765,
  -0.000120789419445943, -0.0173682326446776,
  0.00283358966501266, 0.0189973287452916,
  0.00422780199071588, 0.0190052973194259,
  0.00179133121849407, -0.00491403127579826,
  -0.000225207475048401, -0.0107962067977305,
  -1.74722989377611e-06, -0.00740558095890664,
  -0.0010952915153778, -0.0127869281776265,
  -0.0031126377106639, -0.0164159991897284,
  0.00382568321692876, -0.0139746699789109,
  0.00119362192915543, -0.0108838326480225,
  -0.000918524154543078, -0.00373842537552616,
  -0.00453563160937633, -0.00583244462074028,
  0.00203307718693747, 0.00818465605235041,
  2.41433912589821e-05, 0.00277006105992084,
  -2.4143391259698e-05, 0.0027700610599215,
  0.0003562726813651, -0.0021679180711065,
  2.34920430382964e-05, -0.00438769595812971,
  -0.000172123546682139, -0.00254278760316229,
  0.00076709120349705, -0.000971229887305469,
  0, 0,
  0, 0,
  0, 0,
  -0.000978298976467, 0.000436367489985878,
  -0.00345103764311434, 0.000908266229595611,
  0.00412109125589754, 0.00177690767774896,
  0.00097789242659398, -0.00236487402338126,
  4.78692538101127e-05, -0.000224710065450662,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00276153903543144, -0.00631233885812899,
  0.00389639800366504, -0.0156962556786211,
  4.03280713772066e-05, -0.00473029015254078,
  -9.5046275533288e-05, -0.00555475411881501,
  -0.000130939693550574, -0.00694934258454194,
  0.000216838344254877, -0.0080852613143112,
  -0.000266440785664949, -0.000593899363811934,
  -0.00232961279909512, 0.0127932357712632,
  -0.00366305504496651, 0.0102867433563334,
  0.00270756750379579, 0.00773139847813131,
  -0.000702024761447, 0.0131502159691688,
  -0.000864904726914483, 0.0159004440525603,
  0.00106053319037263, 0.00924917457788288,
  -9.43147583366058e-05, 0.00573742999504523,
  -2.50001627276557e-05, 0.00985209757549987,
  -0.000500909345002226, 0.0137098926105053,
  -0.00236670202191081, 0.0136873218310078,
  0.00351676901116397, -0.00102860536305638,
  0.000649841699541068, 0.00695188374463895,
  0.000533453343925147, 0.00302031875200948,
  -0.000175015488388196, -0.000966023983520969,
  -5.78492841729173e-05, -0.00413180363176857,
  -0.00061646711429136, -0.00831796673958407,
  -0.000770920634429311, -0.0101199018372327,
  -0.00414439054297261, -0.0201582122554649,
  0.00116454257327335, -0.011596813418753,
  7.94265624637976e-05, -0.0117378521857061,
  -5.3693563716093e-05, -0.00954668755381394,
  9.85700799303469e-05, -0.00944264500787351,
  9.40619830076136e-05, -0.00048133436534914,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -2.10630584948613e-05, 9.30744247047421e-05,
  -0.000398652748360631, 0.00454880053911144,
  -0.00104922545344898, 0.0097634308418888,
  -0.0034798668807886, 0.0142923340853669,
  0.00279772394042927, -0.0144594198949242,
  0.00128163427276367, -0.000377110104700984,
  8.40724744396133e-05, 3.09276330203723e-05,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.000703669239415099, 0.000722103841071631,
  -0.00163211946018815, 0.00626189071270788,
  0.0028614915963012, -0.0173936477310725,
  0.00165885716299603, -0.0174973632802502,
  0.000549496243478134, -0.0135073671992543,
  -0.00275665916733126, -0.0134780881342296,
  0.00342871297228792, -0.0184280550834377,
  -0.0028123998206996, -0.0170018555658329,
  0.00206610147627808, -0.0137608758020769,
  -0.000364492777619064, -0.0125356071973395,
  -0.000742732168234484, -0.0134766915129945,
  -0.00334570471414719, -0.00928844761034897,
  0.00113291671113947, -0.00937372515981916,
  -0.000109094980454929, -0.00863877893409049,
  -0.000119546589258648, -0.00925729923002216,
  0.000388223912514851, -0.00485163885279505,
  3.0404114440561e-06, -2.23882511487528e-05,
  0, 0,
  -6.56077040229762e-05, -0.000513738399319896,
  -0.000170435795038834, 0.000716906158798825,
  -0.000341134509486687, 0.00766011667780786,
  -0.000499674489107745, 0.0130278363132486,
  -0.00149723390206193, 0.0188135474021609,
  0.00344764431332289, -0.017138563809207,
  0.00137702810341985, -0.0160255978392951,
  0.000452922888849166, -0.0124685525205037,
  0.000249831937810137, -0.00959732153820858,
  0.000157346664841111, -0.0071011194451911,
  0.000109135951257989, -0.00492630623253532,
  8.73834587981656e-05, -0.00303692506283215,
  6.7879127131063e-05, -0.0013435862623894,
  1.12817628814099e-05, -8.92889767385441e-05,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -2.61984845847785e-05, -0.000219230622539257,
  2.16191772352962e-05, -0.000792288388377083,
  -0.000484194542769407, -0.00667605523635584,
  3.13341471391048e-05, -0.00816943594447528,
  -4.21439882086045e-05, -0.00754424528908526,
  -0.00109024473521979, -0.00948905145163437,
  0.000130863301961551, -0.0169120588084606,
  -0.00232772844100849, -0.019325157515274,
  -0.00268630703788605, -0.0168918072823845,
  0.00164928123611206, -0.0166651437942851,
  0.000228960868256117, -0.0120531548542677,
  -0.000424846547708799, -0.0131102200239654,
  -0.000706007458523082, -0.0152849264820676,
  -0.00263911615585417, -0.011506716399968,
  0.00239916202035495, -0.0187615530271665,
  0.000572195057191347, -0.0155496307733405,
  0.000274924618383192, -0.0139616076547542,
  0.000197559517089947, -0.0128009547096484,
  0.000115931609993653, -0.0116919933568276,
  8.17259176040159e-05, -0.0107944424234607,
  7.88149734088177e-05, -0.0100634934104447,
  -0.00234627269340662, -0.0366266259930517 ;

 tile2_distance =
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _,
  _, _ ;
}
